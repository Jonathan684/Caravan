magic
tech sky130A
magscale 1 2
timestamp 1712065364
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 1104 76 558808 349840
<< metal2 >>
rect 10046 0 10102 800
rect 11150 0 11206 800
rect 12254 0 12310 800
rect 13358 0 13414 800
rect 14462 0 14518 800
rect 15566 0 15622 800
rect 16670 0 16726 800
rect 17774 0 17830 800
rect 18878 0 18934 800
rect 19982 0 20038 800
rect 21086 0 21142 800
rect 22190 0 22246 800
rect 23294 0 23350 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26606 0 26662 800
rect 27710 0 27766 800
rect 28814 0 28870 800
rect 29918 0 29974 800
rect 31022 0 31078 800
rect 32126 0 32182 800
rect 33230 0 33286 800
rect 34334 0 34390 800
rect 35438 0 35494 800
rect 36542 0 36598 800
rect 37646 0 37702 800
rect 38750 0 38806 800
rect 39854 0 39910 800
rect 40958 0 41014 800
rect 42062 0 42118 800
rect 43166 0 43222 800
rect 44270 0 44326 800
rect 45374 0 45430 800
rect 46478 0 46534 800
rect 47582 0 47638 800
rect 48686 0 48742 800
rect 49790 0 49846 800
rect 50894 0 50950 800
rect 51998 0 52054 800
rect 53102 0 53158 800
rect 54206 0 54262 800
rect 55310 0 55366 800
rect 56414 0 56470 800
rect 57518 0 57574 800
rect 58622 0 58678 800
rect 59726 0 59782 800
rect 60830 0 60886 800
rect 61934 0 61990 800
rect 63038 0 63094 800
rect 64142 0 64198 800
rect 65246 0 65302 800
rect 66350 0 66406 800
rect 67454 0 67510 800
rect 68558 0 68614 800
rect 69662 0 69718 800
rect 70766 0 70822 800
rect 71870 0 71926 800
rect 72974 0 73030 800
rect 74078 0 74134 800
rect 75182 0 75238 800
rect 76286 0 76342 800
rect 77390 0 77446 800
rect 78494 0 78550 800
rect 79598 0 79654 800
rect 80702 0 80758 800
rect 81806 0 81862 800
rect 82910 0 82966 800
rect 84014 0 84070 800
rect 85118 0 85174 800
rect 86222 0 86278 800
rect 87326 0 87382 800
rect 88430 0 88486 800
rect 89534 0 89590 800
rect 90638 0 90694 800
rect 91742 0 91798 800
rect 92846 0 92902 800
rect 93950 0 94006 800
rect 95054 0 95110 800
rect 96158 0 96214 800
rect 97262 0 97318 800
rect 98366 0 98422 800
rect 99470 0 99526 800
rect 100574 0 100630 800
rect 101678 0 101734 800
rect 102782 0 102838 800
rect 103886 0 103942 800
rect 104990 0 105046 800
rect 106094 0 106150 800
rect 107198 0 107254 800
rect 108302 0 108358 800
rect 109406 0 109462 800
rect 110510 0 110566 800
rect 111614 0 111670 800
rect 112718 0 112774 800
rect 113822 0 113878 800
rect 114926 0 114982 800
rect 116030 0 116086 800
rect 117134 0 117190 800
rect 118238 0 118294 800
rect 119342 0 119398 800
rect 120446 0 120502 800
rect 121550 0 121606 800
rect 122654 0 122710 800
rect 123758 0 123814 800
rect 124862 0 124918 800
rect 125966 0 126022 800
rect 127070 0 127126 800
rect 128174 0 128230 800
rect 129278 0 129334 800
rect 130382 0 130438 800
rect 131486 0 131542 800
rect 132590 0 132646 800
rect 133694 0 133750 800
rect 134798 0 134854 800
rect 135902 0 135958 800
rect 137006 0 137062 800
rect 138110 0 138166 800
rect 139214 0 139270 800
rect 140318 0 140374 800
rect 141422 0 141478 800
rect 142526 0 142582 800
rect 143630 0 143686 800
rect 144734 0 144790 800
rect 145838 0 145894 800
rect 146942 0 146998 800
rect 148046 0 148102 800
rect 149150 0 149206 800
rect 150254 0 150310 800
rect 151358 0 151414 800
rect 152462 0 152518 800
rect 153566 0 153622 800
rect 154670 0 154726 800
rect 155774 0 155830 800
rect 156878 0 156934 800
rect 157982 0 158038 800
rect 159086 0 159142 800
rect 160190 0 160246 800
rect 161294 0 161350 800
rect 162398 0 162454 800
rect 163502 0 163558 800
rect 164606 0 164662 800
rect 165710 0 165766 800
rect 166814 0 166870 800
rect 167918 0 167974 800
rect 169022 0 169078 800
rect 170126 0 170182 800
rect 171230 0 171286 800
rect 172334 0 172390 800
rect 173438 0 173494 800
rect 174542 0 174598 800
rect 175646 0 175702 800
rect 176750 0 176806 800
rect 177854 0 177910 800
rect 178958 0 179014 800
rect 180062 0 180118 800
rect 181166 0 181222 800
rect 182270 0 182326 800
rect 183374 0 183430 800
rect 184478 0 184534 800
rect 185582 0 185638 800
rect 186686 0 186742 800
rect 187790 0 187846 800
rect 188894 0 188950 800
rect 189998 0 190054 800
rect 191102 0 191158 800
rect 192206 0 192262 800
rect 193310 0 193366 800
rect 194414 0 194470 800
rect 195518 0 195574 800
rect 196622 0 196678 800
rect 197726 0 197782 800
rect 198830 0 198886 800
rect 199934 0 199990 800
rect 201038 0 201094 800
rect 202142 0 202198 800
rect 203246 0 203302 800
rect 204350 0 204406 800
rect 205454 0 205510 800
rect 206558 0 206614 800
rect 207662 0 207718 800
rect 208766 0 208822 800
rect 209870 0 209926 800
rect 210974 0 211030 800
rect 212078 0 212134 800
rect 213182 0 213238 800
rect 214286 0 214342 800
rect 215390 0 215446 800
rect 216494 0 216550 800
rect 217598 0 217654 800
rect 218702 0 218758 800
rect 219806 0 219862 800
rect 220910 0 220966 800
rect 222014 0 222070 800
rect 223118 0 223174 800
rect 224222 0 224278 800
rect 225326 0 225382 800
rect 226430 0 226486 800
rect 227534 0 227590 800
rect 228638 0 228694 800
rect 229742 0 229798 800
rect 230846 0 230902 800
rect 231950 0 232006 800
rect 233054 0 233110 800
rect 234158 0 234214 800
rect 235262 0 235318 800
rect 236366 0 236422 800
rect 237470 0 237526 800
rect 238574 0 238630 800
rect 239678 0 239734 800
rect 240782 0 240838 800
rect 241886 0 241942 800
rect 242990 0 243046 800
rect 244094 0 244150 800
rect 245198 0 245254 800
rect 246302 0 246358 800
rect 247406 0 247462 800
rect 248510 0 248566 800
rect 249614 0 249670 800
rect 250718 0 250774 800
rect 251822 0 251878 800
rect 252926 0 252982 800
rect 254030 0 254086 800
rect 255134 0 255190 800
rect 256238 0 256294 800
rect 257342 0 257398 800
rect 258446 0 258502 800
rect 259550 0 259606 800
rect 260654 0 260710 800
rect 261758 0 261814 800
rect 262862 0 262918 800
rect 263966 0 264022 800
rect 265070 0 265126 800
rect 266174 0 266230 800
rect 267278 0 267334 800
rect 268382 0 268438 800
rect 269486 0 269542 800
rect 270590 0 270646 800
rect 271694 0 271750 800
rect 272798 0 272854 800
rect 273902 0 273958 800
rect 275006 0 275062 800
rect 276110 0 276166 800
rect 277214 0 277270 800
rect 278318 0 278374 800
rect 279422 0 279478 800
rect 280526 0 280582 800
rect 281630 0 281686 800
rect 282734 0 282790 800
rect 283838 0 283894 800
rect 284942 0 284998 800
rect 286046 0 286102 800
rect 287150 0 287206 800
rect 288254 0 288310 800
rect 289358 0 289414 800
rect 290462 0 290518 800
rect 291566 0 291622 800
rect 292670 0 292726 800
rect 293774 0 293830 800
rect 294878 0 294934 800
rect 295982 0 296038 800
rect 297086 0 297142 800
rect 298190 0 298246 800
rect 299294 0 299350 800
rect 300398 0 300454 800
rect 301502 0 301558 800
rect 302606 0 302662 800
rect 303710 0 303766 800
rect 304814 0 304870 800
rect 305918 0 305974 800
rect 307022 0 307078 800
rect 308126 0 308182 800
rect 309230 0 309286 800
rect 310334 0 310390 800
rect 311438 0 311494 800
rect 312542 0 312598 800
rect 313646 0 313702 800
rect 314750 0 314806 800
rect 315854 0 315910 800
rect 316958 0 317014 800
rect 318062 0 318118 800
rect 319166 0 319222 800
rect 320270 0 320326 800
rect 321374 0 321430 800
rect 322478 0 322534 800
rect 323582 0 323638 800
rect 324686 0 324742 800
rect 325790 0 325846 800
rect 326894 0 326950 800
rect 327998 0 328054 800
rect 329102 0 329158 800
rect 330206 0 330262 800
rect 331310 0 331366 800
rect 332414 0 332470 800
rect 333518 0 333574 800
rect 334622 0 334678 800
rect 335726 0 335782 800
rect 336830 0 336886 800
rect 337934 0 337990 800
rect 339038 0 339094 800
rect 340142 0 340198 800
rect 341246 0 341302 800
rect 342350 0 342406 800
rect 343454 0 343510 800
rect 344558 0 344614 800
rect 345662 0 345718 800
rect 346766 0 346822 800
rect 347870 0 347926 800
rect 348974 0 349030 800
rect 350078 0 350134 800
rect 351182 0 351238 800
rect 352286 0 352342 800
rect 353390 0 353446 800
rect 354494 0 354550 800
rect 355598 0 355654 800
rect 356702 0 356758 800
rect 357806 0 357862 800
rect 358910 0 358966 800
rect 360014 0 360070 800
rect 361118 0 361174 800
rect 362222 0 362278 800
rect 363326 0 363382 800
rect 364430 0 364486 800
rect 365534 0 365590 800
rect 366638 0 366694 800
rect 367742 0 367798 800
rect 368846 0 368902 800
rect 369950 0 370006 800
rect 371054 0 371110 800
rect 372158 0 372214 800
rect 373262 0 373318 800
rect 374366 0 374422 800
rect 375470 0 375526 800
rect 376574 0 376630 800
rect 377678 0 377734 800
rect 378782 0 378838 800
rect 379886 0 379942 800
rect 380990 0 381046 800
rect 382094 0 382150 800
rect 383198 0 383254 800
rect 384302 0 384358 800
rect 385406 0 385462 800
rect 386510 0 386566 800
rect 387614 0 387670 800
rect 388718 0 388774 800
rect 389822 0 389878 800
rect 390926 0 390982 800
rect 392030 0 392086 800
rect 393134 0 393190 800
rect 394238 0 394294 800
rect 395342 0 395398 800
rect 396446 0 396502 800
rect 397550 0 397606 800
rect 398654 0 398710 800
rect 399758 0 399814 800
rect 400862 0 400918 800
rect 401966 0 402022 800
rect 403070 0 403126 800
rect 404174 0 404230 800
rect 405278 0 405334 800
rect 406382 0 406438 800
rect 407486 0 407542 800
rect 408590 0 408646 800
rect 409694 0 409750 800
rect 410798 0 410854 800
rect 411902 0 411958 800
rect 413006 0 413062 800
rect 414110 0 414166 800
rect 415214 0 415270 800
rect 416318 0 416374 800
rect 417422 0 417478 800
rect 418526 0 418582 800
rect 419630 0 419686 800
rect 420734 0 420790 800
rect 421838 0 421894 800
rect 422942 0 422998 800
rect 424046 0 424102 800
rect 425150 0 425206 800
rect 426254 0 426310 800
rect 427358 0 427414 800
rect 428462 0 428518 800
rect 429566 0 429622 800
rect 430670 0 430726 800
rect 431774 0 431830 800
rect 432878 0 432934 800
rect 433982 0 434038 800
rect 435086 0 435142 800
rect 436190 0 436246 800
rect 437294 0 437350 800
rect 438398 0 438454 800
rect 439502 0 439558 800
rect 440606 0 440662 800
rect 441710 0 441766 800
rect 442814 0 442870 800
rect 443918 0 443974 800
rect 445022 0 445078 800
rect 446126 0 446182 800
rect 447230 0 447286 800
rect 448334 0 448390 800
rect 449438 0 449494 800
rect 450542 0 450598 800
rect 451646 0 451702 800
rect 452750 0 452806 800
rect 453854 0 453910 800
rect 454958 0 455014 800
rect 456062 0 456118 800
rect 457166 0 457222 800
rect 458270 0 458326 800
rect 459374 0 459430 800
rect 460478 0 460534 800
rect 461582 0 461638 800
rect 462686 0 462742 800
rect 463790 0 463846 800
rect 464894 0 464950 800
rect 465998 0 466054 800
rect 467102 0 467158 800
rect 468206 0 468262 800
rect 469310 0 469366 800
rect 470414 0 470470 800
rect 471518 0 471574 800
rect 472622 0 472678 800
rect 473726 0 473782 800
rect 474830 0 474886 800
rect 475934 0 475990 800
rect 477038 0 477094 800
rect 478142 0 478198 800
rect 479246 0 479302 800
rect 480350 0 480406 800
rect 481454 0 481510 800
rect 482558 0 482614 800
rect 483662 0 483718 800
rect 484766 0 484822 800
rect 485870 0 485926 800
rect 486974 0 487030 800
rect 488078 0 488134 800
rect 489182 0 489238 800
rect 490286 0 490342 800
rect 491390 0 491446 800
rect 492494 0 492550 800
rect 493598 0 493654 800
rect 494702 0 494758 800
rect 495806 0 495862 800
rect 496910 0 496966 800
rect 498014 0 498070 800
rect 499118 0 499174 800
rect 500222 0 500278 800
rect 501326 0 501382 800
rect 502430 0 502486 800
rect 503534 0 503590 800
rect 504638 0 504694 800
rect 505742 0 505798 800
rect 506846 0 506902 800
rect 507950 0 508006 800
rect 509054 0 509110 800
rect 510158 0 510214 800
rect 511262 0 511318 800
rect 512366 0 512422 800
rect 513470 0 513526 800
rect 514574 0 514630 800
rect 515678 0 515734 800
rect 516782 0 516838 800
rect 517886 0 517942 800
rect 518990 0 519046 800
rect 520094 0 520150 800
rect 521198 0 521254 800
rect 522302 0 522358 800
rect 523406 0 523462 800
rect 524510 0 524566 800
rect 525614 0 525670 800
rect 526718 0 526774 800
rect 527822 0 527878 800
rect 528926 0 528982 800
rect 530030 0 530086 800
rect 531134 0 531190 800
rect 532238 0 532294 800
rect 533342 0 533398 800
rect 534446 0 534502 800
rect 535550 0 535606 800
rect 536654 0 536710 800
rect 537758 0 537814 800
rect 538862 0 538918 800
rect 539966 0 540022 800
rect 541070 0 541126 800
rect 542174 0 542230 800
rect 543278 0 543334 800
rect 544382 0 544438 800
rect 545486 0 545542 800
rect 546590 0 546646 800
rect 547694 0 547750 800
rect 548798 0 548854 800
rect 549902 0 549958 800
<< obsm2 >>
rect 1214 856 558420 349829
rect 1214 70 9990 856
rect 10158 70 11094 856
rect 11262 70 12198 856
rect 12366 70 13302 856
rect 13470 70 14406 856
rect 14574 70 15510 856
rect 15678 70 16614 856
rect 16782 70 17718 856
rect 17886 70 18822 856
rect 18990 70 19926 856
rect 20094 70 21030 856
rect 21198 70 22134 856
rect 22302 70 23238 856
rect 23406 70 24342 856
rect 24510 70 25446 856
rect 25614 70 26550 856
rect 26718 70 27654 856
rect 27822 70 28758 856
rect 28926 70 29862 856
rect 30030 70 30966 856
rect 31134 70 32070 856
rect 32238 70 33174 856
rect 33342 70 34278 856
rect 34446 70 35382 856
rect 35550 70 36486 856
rect 36654 70 37590 856
rect 37758 70 38694 856
rect 38862 70 39798 856
rect 39966 70 40902 856
rect 41070 70 42006 856
rect 42174 70 43110 856
rect 43278 70 44214 856
rect 44382 70 45318 856
rect 45486 70 46422 856
rect 46590 70 47526 856
rect 47694 70 48630 856
rect 48798 70 49734 856
rect 49902 70 50838 856
rect 51006 70 51942 856
rect 52110 70 53046 856
rect 53214 70 54150 856
rect 54318 70 55254 856
rect 55422 70 56358 856
rect 56526 70 57462 856
rect 57630 70 58566 856
rect 58734 70 59670 856
rect 59838 70 60774 856
rect 60942 70 61878 856
rect 62046 70 62982 856
rect 63150 70 64086 856
rect 64254 70 65190 856
rect 65358 70 66294 856
rect 66462 70 67398 856
rect 67566 70 68502 856
rect 68670 70 69606 856
rect 69774 70 70710 856
rect 70878 70 71814 856
rect 71982 70 72918 856
rect 73086 70 74022 856
rect 74190 70 75126 856
rect 75294 70 76230 856
rect 76398 70 77334 856
rect 77502 70 78438 856
rect 78606 70 79542 856
rect 79710 70 80646 856
rect 80814 70 81750 856
rect 81918 70 82854 856
rect 83022 70 83958 856
rect 84126 70 85062 856
rect 85230 70 86166 856
rect 86334 70 87270 856
rect 87438 70 88374 856
rect 88542 70 89478 856
rect 89646 70 90582 856
rect 90750 70 91686 856
rect 91854 70 92790 856
rect 92958 70 93894 856
rect 94062 70 94998 856
rect 95166 70 96102 856
rect 96270 70 97206 856
rect 97374 70 98310 856
rect 98478 70 99414 856
rect 99582 70 100518 856
rect 100686 70 101622 856
rect 101790 70 102726 856
rect 102894 70 103830 856
rect 103998 70 104934 856
rect 105102 70 106038 856
rect 106206 70 107142 856
rect 107310 70 108246 856
rect 108414 70 109350 856
rect 109518 70 110454 856
rect 110622 70 111558 856
rect 111726 70 112662 856
rect 112830 70 113766 856
rect 113934 70 114870 856
rect 115038 70 115974 856
rect 116142 70 117078 856
rect 117246 70 118182 856
rect 118350 70 119286 856
rect 119454 70 120390 856
rect 120558 70 121494 856
rect 121662 70 122598 856
rect 122766 70 123702 856
rect 123870 70 124806 856
rect 124974 70 125910 856
rect 126078 70 127014 856
rect 127182 70 128118 856
rect 128286 70 129222 856
rect 129390 70 130326 856
rect 130494 70 131430 856
rect 131598 70 132534 856
rect 132702 70 133638 856
rect 133806 70 134742 856
rect 134910 70 135846 856
rect 136014 70 136950 856
rect 137118 70 138054 856
rect 138222 70 139158 856
rect 139326 70 140262 856
rect 140430 70 141366 856
rect 141534 70 142470 856
rect 142638 70 143574 856
rect 143742 70 144678 856
rect 144846 70 145782 856
rect 145950 70 146886 856
rect 147054 70 147990 856
rect 148158 70 149094 856
rect 149262 70 150198 856
rect 150366 70 151302 856
rect 151470 70 152406 856
rect 152574 70 153510 856
rect 153678 70 154614 856
rect 154782 70 155718 856
rect 155886 70 156822 856
rect 156990 70 157926 856
rect 158094 70 159030 856
rect 159198 70 160134 856
rect 160302 70 161238 856
rect 161406 70 162342 856
rect 162510 70 163446 856
rect 163614 70 164550 856
rect 164718 70 165654 856
rect 165822 70 166758 856
rect 166926 70 167862 856
rect 168030 70 168966 856
rect 169134 70 170070 856
rect 170238 70 171174 856
rect 171342 70 172278 856
rect 172446 70 173382 856
rect 173550 70 174486 856
rect 174654 70 175590 856
rect 175758 70 176694 856
rect 176862 70 177798 856
rect 177966 70 178902 856
rect 179070 70 180006 856
rect 180174 70 181110 856
rect 181278 70 182214 856
rect 182382 70 183318 856
rect 183486 70 184422 856
rect 184590 70 185526 856
rect 185694 70 186630 856
rect 186798 70 187734 856
rect 187902 70 188838 856
rect 189006 70 189942 856
rect 190110 70 191046 856
rect 191214 70 192150 856
rect 192318 70 193254 856
rect 193422 70 194358 856
rect 194526 70 195462 856
rect 195630 70 196566 856
rect 196734 70 197670 856
rect 197838 70 198774 856
rect 198942 70 199878 856
rect 200046 70 200982 856
rect 201150 70 202086 856
rect 202254 70 203190 856
rect 203358 70 204294 856
rect 204462 70 205398 856
rect 205566 70 206502 856
rect 206670 70 207606 856
rect 207774 70 208710 856
rect 208878 70 209814 856
rect 209982 70 210918 856
rect 211086 70 212022 856
rect 212190 70 213126 856
rect 213294 70 214230 856
rect 214398 70 215334 856
rect 215502 70 216438 856
rect 216606 70 217542 856
rect 217710 70 218646 856
rect 218814 70 219750 856
rect 219918 70 220854 856
rect 221022 70 221958 856
rect 222126 70 223062 856
rect 223230 70 224166 856
rect 224334 70 225270 856
rect 225438 70 226374 856
rect 226542 70 227478 856
rect 227646 70 228582 856
rect 228750 70 229686 856
rect 229854 70 230790 856
rect 230958 70 231894 856
rect 232062 70 232998 856
rect 233166 70 234102 856
rect 234270 70 235206 856
rect 235374 70 236310 856
rect 236478 70 237414 856
rect 237582 70 238518 856
rect 238686 70 239622 856
rect 239790 70 240726 856
rect 240894 70 241830 856
rect 241998 70 242934 856
rect 243102 70 244038 856
rect 244206 70 245142 856
rect 245310 70 246246 856
rect 246414 70 247350 856
rect 247518 70 248454 856
rect 248622 70 249558 856
rect 249726 70 250662 856
rect 250830 70 251766 856
rect 251934 70 252870 856
rect 253038 70 253974 856
rect 254142 70 255078 856
rect 255246 70 256182 856
rect 256350 70 257286 856
rect 257454 70 258390 856
rect 258558 70 259494 856
rect 259662 70 260598 856
rect 260766 70 261702 856
rect 261870 70 262806 856
rect 262974 70 263910 856
rect 264078 70 265014 856
rect 265182 70 266118 856
rect 266286 70 267222 856
rect 267390 70 268326 856
rect 268494 70 269430 856
rect 269598 70 270534 856
rect 270702 70 271638 856
rect 271806 70 272742 856
rect 272910 70 273846 856
rect 274014 70 274950 856
rect 275118 70 276054 856
rect 276222 70 277158 856
rect 277326 70 278262 856
rect 278430 70 279366 856
rect 279534 70 280470 856
rect 280638 70 281574 856
rect 281742 70 282678 856
rect 282846 70 283782 856
rect 283950 70 284886 856
rect 285054 70 285990 856
rect 286158 70 287094 856
rect 287262 70 288198 856
rect 288366 70 289302 856
rect 289470 70 290406 856
rect 290574 70 291510 856
rect 291678 70 292614 856
rect 292782 70 293718 856
rect 293886 70 294822 856
rect 294990 70 295926 856
rect 296094 70 297030 856
rect 297198 70 298134 856
rect 298302 70 299238 856
rect 299406 70 300342 856
rect 300510 70 301446 856
rect 301614 70 302550 856
rect 302718 70 303654 856
rect 303822 70 304758 856
rect 304926 70 305862 856
rect 306030 70 306966 856
rect 307134 70 308070 856
rect 308238 70 309174 856
rect 309342 70 310278 856
rect 310446 70 311382 856
rect 311550 70 312486 856
rect 312654 70 313590 856
rect 313758 70 314694 856
rect 314862 70 315798 856
rect 315966 70 316902 856
rect 317070 70 318006 856
rect 318174 70 319110 856
rect 319278 70 320214 856
rect 320382 70 321318 856
rect 321486 70 322422 856
rect 322590 70 323526 856
rect 323694 70 324630 856
rect 324798 70 325734 856
rect 325902 70 326838 856
rect 327006 70 327942 856
rect 328110 70 329046 856
rect 329214 70 330150 856
rect 330318 70 331254 856
rect 331422 70 332358 856
rect 332526 70 333462 856
rect 333630 70 334566 856
rect 334734 70 335670 856
rect 335838 70 336774 856
rect 336942 70 337878 856
rect 338046 70 338982 856
rect 339150 70 340086 856
rect 340254 70 341190 856
rect 341358 70 342294 856
rect 342462 70 343398 856
rect 343566 70 344502 856
rect 344670 70 345606 856
rect 345774 70 346710 856
rect 346878 70 347814 856
rect 347982 70 348918 856
rect 349086 70 350022 856
rect 350190 70 351126 856
rect 351294 70 352230 856
rect 352398 70 353334 856
rect 353502 70 354438 856
rect 354606 70 355542 856
rect 355710 70 356646 856
rect 356814 70 357750 856
rect 357918 70 358854 856
rect 359022 70 359958 856
rect 360126 70 361062 856
rect 361230 70 362166 856
rect 362334 70 363270 856
rect 363438 70 364374 856
rect 364542 70 365478 856
rect 365646 70 366582 856
rect 366750 70 367686 856
rect 367854 70 368790 856
rect 368958 70 369894 856
rect 370062 70 370998 856
rect 371166 70 372102 856
rect 372270 70 373206 856
rect 373374 70 374310 856
rect 374478 70 375414 856
rect 375582 70 376518 856
rect 376686 70 377622 856
rect 377790 70 378726 856
rect 378894 70 379830 856
rect 379998 70 380934 856
rect 381102 70 382038 856
rect 382206 70 383142 856
rect 383310 70 384246 856
rect 384414 70 385350 856
rect 385518 70 386454 856
rect 386622 70 387558 856
rect 387726 70 388662 856
rect 388830 70 389766 856
rect 389934 70 390870 856
rect 391038 70 391974 856
rect 392142 70 393078 856
rect 393246 70 394182 856
rect 394350 70 395286 856
rect 395454 70 396390 856
rect 396558 70 397494 856
rect 397662 70 398598 856
rect 398766 70 399702 856
rect 399870 70 400806 856
rect 400974 70 401910 856
rect 402078 70 403014 856
rect 403182 70 404118 856
rect 404286 70 405222 856
rect 405390 70 406326 856
rect 406494 70 407430 856
rect 407598 70 408534 856
rect 408702 70 409638 856
rect 409806 70 410742 856
rect 410910 70 411846 856
rect 412014 70 412950 856
rect 413118 70 414054 856
rect 414222 70 415158 856
rect 415326 70 416262 856
rect 416430 70 417366 856
rect 417534 70 418470 856
rect 418638 70 419574 856
rect 419742 70 420678 856
rect 420846 70 421782 856
rect 421950 70 422886 856
rect 423054 70 423990 856
rect 424158 70 425094 856
rect 425262 70 426198 856
rect 426366 70 427302 856
rect 427470 70 428406 856
rect 428574 70 429510 856
rect 429678 70 430614 856
rect 430782 70 431718 856
rect 431886 70 432822 856
rect 432990 70 433926 856
rect 434094 70 435030 856
rect 435198 70 436134 856
rect 436302 70 437238 856
rect 437406 70 438342 856
rect 438510 70 439446 856
rect 439614 70 440550 856
rect 440718 70 441654 856
rect 441822 70 442758 856
rect 442926 70 443862 856
rect 444030 70 444966 856
rect 445134 70 446070 856
rect 446238 70 447174 856
rect 447342 70 448278 856
rect 448446 70 449382 856
rect 449550 70 450486 856
rect 450654 70 451590 856
rect 451758 70 452694 856
rect 452862 70 453798 856
rect 453966 70 454902 856
rect 455070 70 456006 856
rect 456174 70 457110 856
rect 457278 70 458214 856
rect 458382 70 459318 856
rect 459486 70 460422 856
rect 460590 70 461526 856
rect 461694 70 462630 856
rect 462798 70 463734 856
rect 463902 70 464838 856
rect 465006 70 465942 856
rect 466110 70 467046 856
rect 467214 70 468150 856
rect 468318 70 469254 856
rect 469422 70 470358 856
rect 470526 70 471462 856
rect 471630 70 472566 856
rect 472734 70 473670 856
rect 473838 70 474774 856
rect 474942 70 475878 856
rect 476046 70 476982 856
rect 477150 70 478086 856
rect 478254 70 479190 856
rect 479358 70 480294 856
rect 480462 70 481398 856
rect 481566 70 482502 856
rect 482670 70 483606 856
rect 483774 70 484710 856
rect 484878 70 485814 856
rect 485982 70 486918 856
rect 487086 70 488022 856
rect 488190 70 489126 856
rect 489294 70 490230 856
rect 490398 70 491334 856
rect 491502 70 492438 856
rect 492606 70 493542 856
rect 493710 70 494646 856
rect 494814 70 495750 856
rect 495918 70 496854 856
rect 497022 70 497958 856
rect 498126 70 499062 856
rect 499230 70 500166 856
rect 500334 70 501270 856
rect 501438 70 502374 856
rect 502542 70 503478 856
rect 503646 70 504582 856
rect 504750 70 505686 856
rect 505854 70 506790 856
rect 506958 70 507894 856
rect 508062 70 508998 856
rect 509166 70 510102 856
rect 510270 70 511206 856
rect 511374 70 512310 856
rect 512478 70 513414 856
rect 513582 70 514518 856
rect 514686 70 515622 856
rect 515790 70 516726 856
rect 516894 70 517830 856
rect 517998 70 518934 856
rect 519102 70 520038 856
rect 520206 70 521142 856
rect 521310 70 522246 856
rect 522414 70 523350 856
rect 523518 70 524454 856
rect 524622 70 525558 856
rect 525726 70 526662 856
rect 526830 70 527766 856
rect 527934 70 528870 856
rect 529038 70 529974 856
rect 530142 70 531078 856
rect 531246 70 532182 856
rect 532350 70 533286 856
rect 533454 70 534390 856
rect 534558 70 535494 856
rect 535662 70 536598 856
rect 536766 70 537702 856
rect 537870 70 538806 856
rect 538974 70 539910 856
rect 540078 70 541014 856
rect 541182 70 542118 856
rect 542286 70 543222 856
rect 543390 70 544326 856
rect 544494 70 545430 856
rect 545598 70 546534 856
rect 546702 70 547638 856
rect 547806 70 548742 856
rect 548910 70 549846 856
rect 550014 70 558420 856
<< metal3 >>
rect 0 341640 800 341760
rect 559200 341640 560000 341760
rect 0 327224 800 327344
rect 559200 327224 560000 327344
rect 0 312808 800 312928
rect 559200 312808 560000 312928
rect 0 298392 800 298512
rect 559200 298392 560000 298512
rect 0 283976 800 284096
rect 559200 283976 560000 284096
rect 0 269560 800 269680
rect 559200 269560 560000 269680
rect 0 255144 800 255264
rect 559200 255144 560000 255264
rect 0 240728 800 240848
rect 559200 240728 560000 240848
rect 0 226312 800 226432
rect 559200 226312 560000 226432
rect 0 211896 800 212016
rect 559200 211896 560000 212016
rect 0 197480 800 197600
rect 559200 197480 560000 197600
rect 0 183064 800 183184
rect 559200 183064 560000 183184
rect 0 168648 800 168768
rect 559200 168648 560000 168768
rect 0 154232 800 154352
rect 559200 154232 560000 154352
rect 0 139816 800 139936
rect 559200 139816 560000 139936
rect 0 125400 800 125520
rect 559200 125400 560000 125520
rect 0 110984 800 111104
rect 559200 110984 560000 111104
rect 0 96568 800 96688
rect 559200 96568 560000 96688
rect 0 82152 800 82272
rect 559200 82152 560000 82272
rect 0 67736 800 67856
rect 559200 67736 560000 67856
rect 0 53320 800 53440
rect 559200 53320 560000 53440
rect 0 38904 800 39024
rect 559200 38904 560000 39024
rect 0 24488 800 24608
rect 559200 24488 560000 24608
rect 0 10072 800 10192
rect 559200 10072 560000 10192
<< obsm3 >>
rect 800 341840 559200 349825
rect 880 341560 559120 341840
rect 800 327424 559200 341560
rect 880 327144 559120 327424
rect 800 313008 559200 327144
rect 880 312728 559120 313008
rect 800 298592 559200 312728
rect 880 298312 559120 298592
rect 800 284176 559200 298312
rect 880 283896 559120 284176
rect 800 269760 559200 283896
rect 880 269480 559120 269760
rect 800 255344 559200 269480
rect 880 255064 559120 255344
rect 800 240928 559200 255064
rect 880 240648 559120 240928
rect 800 226512 559200 240648
rect 880 226232 559120 226512
rect 800 212096 559200 226232
rect 880 211816 559120 212096
rect 800 197680 559200 211816
rect 880 197400 559120 197680
rect 800 183264 559200 197400
rect 880 182984 559120 183264
rect 800 168848 559200 182984
rect 880 168568 559120 168848
rect 800 154432 559200 168568
rect 880 154152 559120 154432
rect 800 140016 559200 154152
rect 880 139736 559120 140016
rect 800 125600 559200 139736
rect 880 125320 559120 125600
rect 800 111184 559200 125320
rect 880 110904 559120 111184
rect 800 96768 559200 110904
rect 880 96488 559120 96768
rect 800 82352 559200 96488
rect 880 82072 559120 82352
rect 800 67936 559200 82072
rect 880 67656 559120 67936
rect 800 53520 559200 67656
rect 880 53240 559120 53520
rect 800 39104 559200 53240
rect 880 38824 559120 39104
rect 800 24688 559200 38824
rect 880 24408 559120 24688
rect 800 10272 559200 24408
rect 880 9992 559120 10272
rect 800 1123 559200 9992
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< obsm4 >>
rect 260603 3979 265248 7173
rect 265728 3979 266005 7173
<< labels >>
rlabel metal3 s 559200 10072 560000 10192 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 255144 800 255264 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 211896 800 212016 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 168648 800 168768 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 559200 53320 560000 53440 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 559200 96568 560000 96688 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 559200 139816 560000 139936 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 559200 183064 560000 183184 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 559200 226312 560000 226432 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 559200 269560 560000 269680 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 559200 312808 560000 312928 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 341640 800 341760 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 298392 800 298512 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 559200 38904 560000 39024 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 226312 800 226432 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 183064 800 183184 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 559200 82152 560000 82272 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 559200 125400 560000 125520 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 559200 168648 560000 168768 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 559200 211896 560000 212016 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 559200 255144 560000 255264 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 559200 298392 560000 298512 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 559200 341640 560000 341760 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 312808 800 312928 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 269560 800 269680 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 559200 24488 560000 24608 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 240728 800 240848 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 197480 800 197600 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 154232 800 154352 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 559200 67736 560000 67856 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 559200 110984 560000 111104 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 559200 154232 560000 154352 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 559200 197480 560000 197600 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 559200 240728 560000 240848 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 559200 283976 560000 284096 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 559200 327224 560000 327344 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 327224 800 327344 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 283976 800 284096 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_in[0]
port 49 nsew signal input
rlabel metal2 s 458270 0 458326 800 6 la_data_in[100]
port 50 nsew signal input
rlabel metal2 s 461582 0 461638 800 6 la_data_in[101]
port 51 nsew signal input
rlabel metal2 s 464894 0 464950 800 6 la_data_in[102]
port 52 nsew signal input
rlabel metal2 s 468206 0 468262 800 6 la_data_in[103]
port 53 nsew signal input
rlabel metal2 s 471518 0 471574 800 6 la_data_in[104]
port 54 nsew signal input
rlabel metal2 s 474830 0 474886 800 6 la_data_in[105]
port 55 nsew signal input
rlabel metal2 s 478142 0 478198 800 6 la_data_in[106]
port 56 nsew signal input
rlabel metal2 s 481454 0 481510 800 6 la_data_in[107]
port 57 nsew signal input
rlabel metal2 s 484766 0 484822 800 6 la_data_in[108]
port 58 nsew signal input
rlabel metal2 s 488078 0 488134 800 6 la_data_in[109]
port 59 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_data_in[10]
port 60 nsew signal input
rlabel metal2 s 491390 0 491446 800 6 la_data_in[110]
port 61 nsew signal input
rlabel metal2 s 494702 0 494758 800 6 la_data_in[111]
port 62 nsew signal input
rlabel metal2 s 498014 0 498070 800 6 la_data_in[112]
port 63 nsew signal input
rlabel metal2 s 501326 0 501382 800 6 la_data_in[113]
port 64 nsew signal input
rlabel metal2 s 504638 0 504694 800 6 la_data_in[114]
port 65 nsew signal input
rlabel metal2 s 507950 0 508006 800 6 la_data_in[115]
port 66 nsew signal input
rlabel metal2 s 511262 0 511318 800 6 la_data_in[116]
port 67 nsew signal input
rlabel metal2 s 514574 0 514630 800 6 la_data_in[117]
port 68 nsew signal input
rlabel metal2 s 517886 0 517942 800 6 la_data_in[118]
port 69 nsew signal input
rlabel metal2 s 521198 0 521254 800 6 la_data_in[119]
port 70 nsew signal input
rlabel metal2 s 163502 0 163558 800 6 la_data_in[11]
port 71 nsew signal input
rlabel metal2 s 524510 0 524566 800 6 la_data_in[120]
port 72 nsew signal input
rlabel metal2 s 527822 0 527878 800 6 la_data_in[121]
port 73 nsew signal input
rlabel metal2 s 531134 0 531190 800 6 la_data_in[122]
port 74 nsew signal input
rlabel metal2 s 534446 0 534502 800 6 la_data_in[123]
port 75 nsew signal input
rlabel metal2 s 537758 0 537814 800 6 la_data_in[124]
port 76 nsew signal input
rlabel metal2 s 541070 0 541126 800 6 la_data_in[125]
port 77 nsew signal input
rlabel metal2 s 544382 0 544438 800 6 la_data_in[126]
port 78 nsew signal input
rlabel metal2 s 547694 0 547750 800 6 la_data_in[127]
port 79 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_data_in[12]
port 80 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_data_in[13]
port 81 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 la_data_in[14]
port 82 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_data_in[15]
port 83 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_data_in[16]
port 84 nsew signal input
rlabel metal2 s 183374 0 183430 800 6 la_data_in[17]
port 85 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 la_data_in[18]
port 86 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_data_in[19]
port 87 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[1]
port 88 nsew signal input
rlabel metal2 s 193310 0 193366 800 6 la_data_in[20]
port 89 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 la_data_in[21]
port 90 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_data_in[22]
port 91 nsew signal input
rlabel metal2 s 203246 0 203302 800 6 la_data_in[23]
port 92 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_data_in[24]
port 93 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_data_in[25]
port 94 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_data_in[26]
port 95 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_data_in[27]
port 96 nsew signal input
rlabel metal2 s 219806 0 219862 800 6 la_data_in[28]
port 97 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_data_in[29]
port 98 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_data_in[2]
port 99 nsew signal input
rlabel metal2 s 226430 0 226486 800 6 la_data_in[30]
port 100 nsew signal input
rlabel metal2 s 229742 0 229798 800 6 la_data_in[31]
port 101 nsew signal input
rlabel metal2 s 233054 0 233110 800 6 la_data_in[32]
port 102 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_data_in[33]
port 103 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_data_in[34]
port 104 nsew signal input
rlabel metal2 s 242990 0 243046 800 6 la_data_in[35]
port 105 nsew signal input
rlabel metal2 s 246302 0 246358 800 6 la_data_in[36]
port 106 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 la_data_in[37]
port 107 nsew signal input
rlabel metal2 s 252926 0 252982 800 6 la_data_in[38]
port 108 nsew signal input
rlabel metal2 s 256238 0 256294 800 6 la_data_in[39]
port 109 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_data_in[3]
port 110 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_data_in[40]
port 111 nsew signal input
rlabel metal2 s 262862 0 262918 800 6 la_data_in[41]
port 112 nsew signal input
rlabel metal2 s 266174 0 266230 800 6 la_data_in[42]
port 113 nsew signal input
rlabel metal2 s 269486 0 269542 800 6 la_data_in[43]
port 114 nsew signal input
rlabel metal2 s 272798 0 272854 800 6 la_data_in[44]
port 115 nsew signal input
rlabel metal2 s 276110 0 276166 800 6 la_data_in[45]
port 116 nsew signal input
rlabel metal2 s 279422 0 279478 800 6 la_data_in[46]
port 117 nsew signal input
rlabel metal2 s 282734 0 282790 800 6 la_data_in[47]
port 118 nsew signal input
rlabel metal2 s 286046 0 286102 800 6 la_data_in[48]
port 119 nsew signal input
rlabel metal2 s 289358 0 289414 800 6 la_data_in[49]
port 120 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_data_in[4]
port 121 nsew signal input
rlabel metal2 s 292670 0 292726 800 6 la_data_in[50]
port 122 nsew signal input
rlabel metal2 s 295982 0 296038 800 6 la_data_in[51]
port 123 nsew signal input
rlabel metal2 s 299294 0 299350 800 6 la_data_in[52]
port 124 nsew signal input
rlabel metal2 s 302606 0 302662 800 6 la_data_in[53]
port 125 nsew signal input
rlabel metal2 s 305918 0 305974 800 6 la_data_in[54]
port 126 nsew signal input
rlabel metal2 s 309230 0 309286 800 6 la_data_in[55]
port 127 nsew signal input
rlabel metal2 s 312542 0 312598 800 6 la_data_in[56]
port 128 nsew signal input
rlabel metal2 s 315854 0 315910 800 6 la_data_in[57]
port 129 nsew signal input
rlabel metal2 s 319166 0 319222 800 6 la_data_in[58]
port 130 nsew signal input
rlabel metal2 s 322478 0 322534 800 6 la_data_in[59]
port 131 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_data_in[5]
port 132 nsew signal input
rlabel metal2 s 325790 0 325846 800 6 la_data_in[60]
port 133 nsew signal input
rlabel metal2 s 329102 0 329158 800 6 la_data_in[61]
port 134 nsew signal input
rlabel metal2 s 332414 0 332470 800 6 la_data_in[62]
port 135 nsew signal input
rlabel metal2 s 335726 0 335782 800 6 la_data_in[63]
port 136 nsew signal input
rlabel metal2 s 339038 0 339094 800 6 la_data_in[64]
port 137 nsew signal input
rlabel metal2 s 342350 0 342406 800 6 la_data_in[65]
port 138 nsew signal input
rlabel metal2 s 345662 0 345718 800 6 la_data_in[66]
port 139 nsew signal input
rlabel metal2 s 348974 0 349030 800 6 la_data_in[67]
port 140 nsew signal input
rlabel metal2 s 352286 0 352342 800 6 la_data_in[68]
port 141 nsew signal input
rlabel metal2 s 355598 0 355654 800 6 la_data_in[69]
port 142 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_data_in[6]
port 143 nsew signal input
rlabel metal2 s 358910 0 358966 800 6 la_data_in[70]
port 144 nsew signal input
rlabel metal2 s 362222 0 362278 800 6 la_data_in[71]
port 145 nsew signal input
rlabel metal2 s 365534 0 365590 800 6 la_data_in[72]
port 146 nsew signal input
rlabel metal2 s 368846 0 368902 800 6 la_data_in[73]
port 147 nsew signal input
rlabel metal2 s 372158 0 372214 800 6 la_data_in[74]
port 148 nsew signal input
rlabel metal2 s 375470 0 375526 800 6 la_data_in[75]
port 149 nsew signal input
rlabel metal2 s 378782 0 378838 800 6 la_data_in[76]
port 150 nsew signal input
rlabel metal2 s 382094 0 382150 800 6 la_data_in[77]
port 151 nsew signal input
rlabel metal2 s 385406 0 385462 800 6 la_data_in[78]
port 152 nsew signal input
rlabel metal2 s 388718 0 388774 800 6 la_data_in[79]
port 153 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_data_in[7]
port 154 nsew signal input
rlabel metal2 s 392030 0 392086 800 6 la_data_in[80]
port 155 nsew signal input
rlabel metal2 s 395342 0 395398 800 6 la_data_in[81]
port 156 nsew signal input
rlabel metal2 s 398654 0 398710 800 6 la_data_in[82]
port 157 nsew signal input
rlabel metal2 s 401966 0 402022 800 6 la_data_in[83]
port 158 nsew signal input
rlabel metal2 s 405278 0 405334 800 6 la_data_in[84]
port 159 nsew signal input
rlabel metal2 s 408590 0 408646 800 6 la_data_in[85]
port 160 nsew signal input
rlabel metal2 s 411902 0 411958 800 6 la_data_in[86]
port 161 nsew signal input
rlabel metal2 s 415214 0 415270 800 6 la_data_in[87]
port 162 nsew signal input
rlabel metal2 s 418526 0 418582 800 6 la_data_in[88]
port 163 nsew signal input
rlabel metal2 s 421838 0 421894 800 6 la_data_in[89]
port 164 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_data_in[8]
port 165 nsew signal input
rlabel metal2 s 425150 0 425206 800 6 la_data_in[90]
port 166 nsew signal input
rlabel metal2 s 428462 0 428518 800 6 la_data_in[91]
port 167 nsew signal input
rlabel metal2 s 431774 0 431830 800 6 la_data_in[92]
port 168 nsew signal input
rlabel metal2 s 435086 0 435142 800 6 la_data_in[93]
port 169 nsew signal input
rlabel metal2 s 438398 0 438454 800 6 la_data_in[94]
port 170 nsew signal input
rlabel metal2 s 441710 0 441766 800 6 la_data_in[95]
port 171 nsew signal input
rlabel metal2 s 445022 0 445078 800 6 la_data_in[96]
port 172 nsew signal input
rlabel metal2 s 448334 0 448390 800 6 la_data_in[97]
port 173 nsew signal input
rlabel metal2 s 451646 0 451702 800 6 la_data_in[98]
port 174 nsew signal input
rlabel metal2 s 454958 0 455014 800 6 la_data_in[99]
port 175 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_data_in[9]
port 176 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_data_out[0]
port 177 nsew signal output
rlabel metal2 s 459374 0 459430 800 6 la_data_out[100]
port 178 nsew signal output
rlabel metal2 s 462686 0 462742 800 6 la_data_out[101]
port 179 nsew signal output
rlabel metal2 s 465998 0 466054 800 6 la_data_out[102]
port 180 nsew signal output
rlabel metal2 s 469310 0 469366 800 6 la_data_out[103]
port 181 nsew signal output
rlabel metal2 s 472622 0 472678 800 6 la_data_out[104]
port 182 nsew signal output
rlabel metal2 s 475934 0 475990 800 6 la_data_out[105]
port 183 nsew signal output
rlabel metal2 s 479246 0 479302 800 6 la_data_out[106]
port 184 nsew signal output
rlabel metal2 s 482558 0 482614 800 6 la_data_out[107]
port 185 nsew signal output
rlabel metal2 s 485870 0 485926 800 6 la_data_out[108]
port 186 nsew signal output
rlabel metal2 s 489182 0 489238 800 6 la_data_out[109]
port 187 nsew signal output
rlabel metal2 s 161294 0 161350 800 6 la_data_out[10]
port 188 nsew signal output
rlabel metal2 s 492494 0 492550 800 6 la_data_out[110]
port 189 nsew signal output
rlabel metal2 s 495806 0 495862 800 6 la_data_out[111]
port 190 nsew signal output
rlabel metal2 s 499118 0 499174 800 6 la_data_out[112]
port 191 nsew signal output
rlabel metal2 s 502430 0 502486 800 6 la_data_out[113]
port 192 nsew signal output
rlabel metal2 s 505742 0 505798 800 6 la_data_out[114]
port 193 nsew signal output
rlabel metal2 s 509054 0 509110 800 6 la_data_out[115]
port 194 nsew signal output
rlabel metal2 s 512366 0 512422 800 6 la_data_out[116]
port 195 nsew signal output
rlabel metal2 s 515678 0 515734 800 6 la_data_out[117]
port 196 nsew signal output
rlabel metal2 s 518990 0 519046 800 6 la_data_out[118]
port 197 nsew signal output
rlabel metal2 s 522302 0 522358 800 6 la_data_out[119]
port 198 nsew signal output
rlabel metal2 s 164606 0 164662 800 6 la_data_out[11]
port 199 nsew signal output
rlabel metal2 s 525614 0 525670 800 6 la_data_out[120]
port 200 nsew signal output
rlabel metal2 s 528926 0 528982 800 6 la_data_out[121]
port 201 nsew signal output
rlabel metal2 s 532238 0 532294 800 6 la_data_out[122]
port 202 nsew signal output
rlabel metal2 s 535550 0 535606 800 6 la_data_out[123]
port 203 nsew signal output
rlabel metal2 s 538862 0 538918 800 6 la_data_out[124]
port 204 nsew signal output
rlabel metal2 s 542174 0 542230 800 6 la_data_out[125]
port 205 nsew signal output
rlabel metal2 s 545486 0 545542 800 6 la_data_out[126]
port 206 nsew signal output
rlabel metal2 s 548798 0 548854 800 6 la_data_out[127]
port 207 nsew signal output
rlabel metal2 s 167918 0 167974 800 6 la_data_out[12]
port 208 nsew signal output
rlabel metal2 s 171230 0 171286 800 6 la_data_out[13]
port 209 nsew signal output
rlabel metal2 s 174542 0 174598 800 6 la_data_out[14]
port 210 nsew signal output
rlabel metal2 s 177854 0 177910 800 6 la_data_out[15]
port 211 nsew signal output
rlabel metal2 s 181166 0 181222 800 6 la_data_out[16]
port 212 nsew signal output
rlabel metal2 s 184478 0 184534 800 6 la_data_out[17]
port 213 nsew signal output
rlabel metal2 s 187790 0 187846 800 6 la_data_out[18]
port 214 nsew signal output
rlabel metal2 s 191102 0 191158 800 6 la_data_out[19]
port 215 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[1]
port 216 nsew signal output
rlabel metal2 s 194414 0 194470 800 6 la_data_out[20]
port 217 nsew signal output
rlabel metal2 s 197726 0 197782 800 6 la_data_out[21]
port 218 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 la_data_out[22]
port 219 nsew signal output
rlabel metal2 s 204350 0 204406 800 6 la_data_out[23]
port 220 nsew signal output
rlabel metal2 s 207662 0 207718 800 6 la_data_out[24]
port 221 nsew signal output
rlabel metal2 s 210974 0 211030 800 6 la_data_out[25]
port 222 nsew signal output
rlabel metal2 s 214286 0 214342 800 6 la_data_out[26]
port 223 nsew signal output
rlabel metal2 s 217598 0 217654 800 6 la_data_out[27]
port 224 nsew signal output
rlabel metal2 s 220910 0 220966 800 6 la_data_out[28]
port 225 nsew signal output
rlabel metal2 s 224222 0 224278 800 6 la_data_out[29]
port 226 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[2]
port 227 nsew signal output
rlabel metal2 s 227534 0 227590 800 6 la_data_out[30]
port 228 nsew signal output
rlabel metal2 s 230846 0 230902 800 6 la_data_out[31]
port 229 nsew signal output
rlabel metal2 s 234158 0 234214 800 6 la_data_out[32]
port 230 nsew signal output
rlabel metal2 s 237470 0 237526 800 6 la_data_out[33]
port 231 nsew signal output
rlabel metal2 s 240782 0 240838 800 6 la_data_out[34]
port 232 nsew signal output
rlabel metal2 s 244094 0 244150 800 6 la_data_out[35]
port 233 nsew signal output
rlabel metal2 s 247406 0 247462 800 6 la_data_out[36]
port 234 nsew signal output
rlabel metal2 s 250718 0 250774 800 6 la_data_out[37]
port 235 nsew signal output
rlabel metal2 s 254030 0 254086 800 6 la_data_out[38]
port 236 nsew signal output
rlabel metal2 s 257342 0 257398 800 6 la_data_out[39]
port 237 nsew signal output
rlabel metal2 s 138110 0 138166 800 6 la_data_out[3]
port 238 nsew signal output
rlabel metal2 s 260654 0 260710 800 6 la_data_out[40]
port 239 nsew signal output
rlabel metal2 s 263966 0 264022 800 6 la_data_out[41]
port 240 nsew signal output
rlabel metal2 s 267278 0 267334 800 6 la_data_out[42]
port 241 nsew signal output
rlabel metal2 s 270590 0 270646 800 6 la_data_out[43]
port 242 nsew signal output
rlabel metal2 s 273902 0 273958 800 6 la_data_out[44]
port 243 nsew signal output
rlabel metal2 s 277214 0 277270 800 6 la_data_out[45]
port 244 nsew signal output
rlabel metal2 s 280526 0 280582 800 6 la_data_out[46]
port 245 nsew signal output
rlabel metal2 s 283838 0 283894 800 6 la_data_out[47]
port 246 nsew signal output
rlabel metal2 s 287150 0 287206 800 6 la_data_out[48]
port 247 nsew signal output
rlabel metal2 s 290462 0 290518 800 6 la_data_out[49]
port 248 nsew signal output
rlabel metal2 s 141422 0 141478 800 6 la_data_out[4]
port 249 nsew signal output
rlabel metal2 s 293774 0 293830 800 6 la_data_out[50]
port 250 nsew signal output
rlabel metal2 s 297086 0 297142 800 6 la_data_out[51]
port 251 nsew signal output
rlabel metal2 s 300398 0 300454 800 6 la_data_out[52]
port 252 nsew signal output
rlabel metal2 s 303710 0 303766 800 6 la_data_out[53]
port 253 nsew signal output
rlabel metal2 s 307022 0 307078 800 6 la_data_out[54]
port 254 nsew signal output
rlabel metal2 s 310334 0 310390 800 6 la_data_out[55]
port 255 nsew signal output
rlabel metal2 s 313646 0 313702 800 6 la_data_out[56]
port 256 nsew signal output
rlabel metal2 s 316958 0 317014 800 6 la_data_out[57]
port 257 nsew signal output
rlabel metal2 s 320270 0 320326 800 6 la_data_out[58]
port 258 nsew signal output
rlabel metal2 s 323582 0 323638 800 6 la_data_out[59]
port 259 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 la_data_out[5]
port 260 nsew signal output
rlabel metal2 s 326894 0 326950 800 6 la_data_out[60]
port 261 nsew signal output
rlabel metal2 s 330206 0 330262 800 6 la_data_out[61]
port 262 nsew signal output
rlabel metal2 s 333518 0 333574 800 6 la_data_out[62]
port 263 nsew signal output
rlabel metal2 s 336830 0 336886 800 6 la_data_out[63]
port 264 nsew signal output
rlabel metal2 s 340142 0 340198 800 6 la_data_out[64]
port 265 nsew signal output
rlabel metal2 s 343454 0 343510 800 6 la_data_out[65]
port 266 nsew signal output
rlabel metal2 s 346766 0 346822 800 6 la_data_out[66]
port 267 nsew signal output
rlabel metal2 s 350078 0 350134 800 6 la_data_out[67]
port 268 nsew signal output
rlabel metal2 s 353390 0 353446 800 6 la_data_out[68]
port 269 nsew signal output
rlabel metal2 s 356702 0 356758 800 6 la_data_out[69]
port 270 nsew signal output
rlabel metal2 s 148046 0 148102 800 6 la_data_out[6]
port 271 nsew signal output
rlabel metal2 s 360014 0 360070 800 6 la_data_out[70]
port 272 nsew signal output
rlabel metal2 s 363326 0 363382 800 6 la_data_out[71]
port 273 nsew signal output
rlabel metal2 s 366638 0 366694 800 6 la_data_out[72]
port 274 nsew signal output
rlabel metal2 s 369950 0 370006 800 6 la_data_out[73]
port 275 nsew signal output
rlabel metal2 s 373262 0 373318 800 6 la_data_out[74]
port 276 nsew signal output
rlabel metal2 s 376574 0 376630 800 6 la_data_out[75]
port 277 nsew signal output
rlabel metal2 s 379886 0 379942 800 6 la_data_out[76]
port 278 nsew signal output
rlabel metal2 s 383198 0 383254 800 6 la_data_out[77]
port 279 nsew signal output
rlabel metal2 s 386510 0 386566 800 6 la_data_out[78]
port 280 nsew signal output
rlabel metal2 s 389822 0 389878 800 6 la_data_out[79]
port 281 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 la_data_out[7]
port 282 nsew signal output
rlabel metal2 s 393134 0 393190 800 6 la_data_out[80]
port 283 nsew signal output
rlabel metal2 s 396446 0 396502 800 6 la_data_out[81]
port 284 nsew signal output
rlabel metal2 s 399758 0 399814 800 6 la_data_out[82]
port 285 nsew signal output
rlabel metal2 s 403070 0 403126 800 6 la_data_out[83]
port 286 nsew signal output
rlabel metal2 s 406382 0 406438 800 6 la_data_out[84]
port 287 nsew signal output
rlabel metal2 s 409694 0 409750 800 6 la_data_out[85]
port 288 nsew signal output
rlabel metal2 s 413006 0 413062 800 6 la_data_out[86]
port 289 nsew signal output
rlabel metal2 s 416318 0 416374 800 6 la_data_out[87]
port 290 nsew signal output
rlabel metal2 s 419630 0 419686 800 6 la_data_out[88]
port 291 nsew signal output
rlabel metal2 s 422942 0 422998 800 6 la_data_out[89]
port 292 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 la_data_out[8]
port 293 nsew signal output
rlabel metal2 s 426254 0 426310 800 6 la_data_out[90]
port 294 nsew signal output
rlabel metal2 s 429566 0 429622 800 6 la_data_out[91]
port 295 nsew signal output
rlabel metal2 s 432878 0 432934 800 6 la_data_out[92]
port 296 nsew signal output
rlabel metal2 s 436190 0 436246 800 6 la_data_out[93]
port 297 nsew signal output
rlabel metal2 s 439502 0 439558 800 6 la_data_out[94]
port 298 nsew signal output
rlabel metal2 s 442814 0 442870 800 6 la_data_out[95]
port 299 nsew signal output
rlabel metal2 s 446126 0 446182 800 6 la_data_out[96]
port 300 nsew signal output
rlabel metal2 s 449438 0 449494 800 6 la_data_out[97]
port 301 nsew signal output
rlabel metal2 s 452750 0 452806 800 6 la_data_out[98]
port 302 nsew signal output
rlabel metal2 s 456062 0 456118 800 6 la_data_out[99]
port 303 nsew signal output
rlabel metal2 s 157982 0 158038 800 6 la_data_out[9]
port 304 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_oenb[0]
port 305 nsew signal input
rlabel metal2 s 460478 0 460534 800 6 la_oenb[100]
port 306 nsew signal input
rlabel metal2 s 463790 0 463846 800 6 la_oenb[101]
port 307 nsew signal input
rlabel metal2 s 467102 0 467158 800 6 la_oenb[102]
port 308 nsew signal input
rlabel metal2 s 470414 0 470470 800 6 la_oenb[103]
port 309 nsew signal input
rlabel metal2 s 473726 0 473782 800 6 la_oenb[104]
port 310 nsew signal input
rlabel metal2 s 477038 0 477094 800 6 la_oenb[105]
port 311 nsew signal input
rlabel metal2 s 480350 0 480406 800 6 la_oenb[106]
port 312 nsew signal input
rlabel metal2 s 483662 0 483718 800 6 la_oenb[107]
port 313 nsew signal input
rlabel metal2 s 486974 0 487030 800 6 la_oenb[108]
port 314 nsew signal input
rlabel metal2 s 490286 0 490342 800 6 la_oenb[109]
port 315 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_oenb[10]
port 316 nsew signal input
rlabel metal2 s 493598 0 493654 800 6 la_oenb[110]
port 317 nsew signal input
rlabel metal2 s 496910 0 496966 800 6 la_oenb[111]
port 318 nsew signal input
rlabel metal2 s 500222 0 500278 800 6 la_oenb[112]
port 319 nsew signal input
rlabel metal2 s 503534 0 503590 800 6 la_oenb[113]
port 320 nsew signal input
rlabel metal2 s 506846 0 506902 800 6 la_oenb[114]
port 321 nsew signal input
rlabel metal2 s 510158 0 510214 800 6 la_oenb[115]
port 322 nsew signal input
rlabel metal2 s 513470 0 513526 800 6 la_oenb[116]
port 323 nsew signal input
rlabel metal2 s 516782 0 516838 800 6 la_oenb[117]
port 324 nsew signal input
rlabel metal2 s 520094 0 520150 800 6 la_oenb[118]
port 325 nsew signal input
rlabel metal2 s 523406 0 523462 800 6 la_oenb[119]
port 326 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_oenb[11]
port 327 nsew signal input
rlabel metal2 s 526718 0 526774 800 6 la_oenb[120]
port 328 nsew signal input
rlabel metal2 s 530030 0 530086 800 6 la_oenb[121]
port 329 nsew signal input
rlabel metal2 s 533342 0 533398 800 6 la_oenb[122]
port 330 nsew signal input
rlabel metal2 s 536654 0 536710 800 6 la_oenb[123]
port 331 nsew signal input
rlabel metal2 s 539966 0 540022 800 6 la_oenb[124]
port 332 nsew signal input
rlabel metal2 s 543278 0 543334 800 6 la_oenb[125]
port 333 nsew signal input
rlabel metal2 s 546590 0 546646 800 6 la_oenb[126]
port 334 nsew signal input
rlabel metal2 s 549902 0 549958 800 6 la_oenb[127]
port 335 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_oenb[12]
port 336 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 la_oenb[13]
port 337 nsew signal input
rlabel metal2 s 175646 0 175702 800 6 la_oenb[14]
port 338 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 la_oenb[15]
port 339 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_oenb[16]
port 340 nsew signal input
rlabel metal2 s 185582 0 185638 800 6 la_oenb[17]
port 341 nsew signal input
rlabel metal2 s 188894 0 188950 800 6 la_oenb[18]
port 342 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 la_oenb[19]
port 343 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_oenb[1]
port 344 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 la_oenb[20]
port 345 nsew signal input
rlabel metal2 s 198830 0 198886 800 6 la_oenb[21]
port 346 nsew signal input
rlabel metal2 s 202142 0 202198 800 6 la_oenb[22]
port 347 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_oenb[23]
port 348 nsew signal input
rlabel metal2 s 208766 0 208822 800 6 la_oenb[24]
port 349 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 la_oenb[25]
port 350 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_oenb[26]
port 351 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_oenb[27]
port 352 nsew signal input
rlabel metal2 s 222014 0 222070 800 6 la_oenb[28]
port 353 nsew signal input
rlabel metal2 s 225326 0 225382 800 6 la_oenb[29]
port 354 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[2]
port 355 nsew signal input
rlabel metal2 s 228638 0 228694 800 6 la_oenb[30]
port 356 nsew signal input
rlabel metal2 s 231950 0 232006 800 6 la_oenb[31]
port 357 nsew signal input
rlabel metal2 s 235262 0 235318 800 6 la_oenb[32]
port 358 nsew signal input
rlabel metal2 s 238574 0 238630 800 6 la_oenb[33]
port 359 nsew signal input
rlabel metal2 s 241886 0 241942 800 6 la_oenb[34]
port 360 nsew signal input
rlabel metal2 s 245198 0 245254 800 6 la_oenb[35]
port 361 nsew signal input
rlabel metal2 s 248510 0 248566 800 6 la_oenb[36]
port 362 nsew signal input
rlabel metal2 s 251822 0 251878 800 6 la_oenb[37]
port 363 nsew signal input
rlabel metal2 s 255134 0 255190 800 6 la_oenb[38]
port 364 nsew signal input
rlabel metal2 s 258446 0 258502 800 6 la_oenb[39]
port 365 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oenb[3]
port 366 nsew signal input
rlabel metal2 s 261758 0 261814 800 6 la_oenb[40]
port 367 nsew signal input
rlabel metal2 s 265070 0 265126 800 6 la_oenb[41]
port 368 nsew signal input
rlabel metal2 s 268382 0 268438 800 6 la_oenb[42]
port 369 nsew signal input
rlabel metal2 s 271694 0 271750 800 6 la_oenb[43]
port 370 nsew signal input
rlabel metal2 s 275006 0 275062 800 6 la_oenb[44]
port 371 nsew signal input
rlabel metal2 s 278318 0 278374 800 6 la_oenb[45]
port 372 nsew signal input
rlabel metal2 s 281630 0 281686 800 6 la_oenb[46]
port 373 nsew signal input
rlabel metal2 s 284942 0 284998 800 6 la_oenb[47]
port 374 nsew signal input
rlabel metal2 s 288254 0 288310 800 6 la_oenb[48]
port 375 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 la_oenb[49]
port 376 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_oenb[4]
port 377 nsew signal input
rlabel metal2 s 294878 0 294934 800 6 la_oenb[50]
port 378 nsew signal input
rlabel metal2 s 298190 0 298246 800 6 la_oenb[51]
port 379 nsew signal input
rlabel metal2 s 301502 0 301558 800 6 la_oenb[52]
port 380 nsew signal input
rlabel metal2 s 304814 0 304870 800 6 la_oenb[53]
port 381 nsew signal input
rlabel metal2 s 308126 0 308182 800 6 la_oenb[54]
port 382 nsew signal input
rlabel metal2 s 311438 0 311494 800 6 la_oenb[55]
port 383 nsew signal input
rlabel metal2 s 314750 0 314806 800 6 la_oenb[56]
port 384 nsew signal input
rlabel metal2 s 318062 0 318118 800 6 la_oenb[57]
port 385 nsew signal input
rlabel metal2 s 321374 0 321430 800 6 la_oenb[58]
port 386 nsew signal input
rlabel metal2 s 324686 0 324742 800 6 la_oenb[59]
port 387 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[5]
port 388 nsew signal input
rlabel metal2 s 327998 0 328054 800 6 la_oenb[60]
port 389 nsew signal input
rlabel metal2 s 331310 0 331366 800 6 la_oenb[61]
port 390 nsew signal input
rlabel metal2 s 334622 0 334678 800 6 la_oenb[62]
port 391 nsew signal input
rlabel metal2 s 337934 0 337990 800 6 la_oenb[63]
port 392 nsew signal input
rlabel metal2 s 341246 0 341302 800 6 la_oenb[64]
port 393 nsew signal input
rlabel metal2 s 344558 0 344614 800 6 la_oenb[65]
port 394 nsew signal input
rlabel metal2 s 347870 0 347926 800 6 la_oenb[66]
port 395 nsew signal input
rlabel metal2 s 351182 0 351238 800 6 la_oenb[67]
port 396 nsew signal input
rlabel metal2 s 354494 0 354550 800 6 la_oenb[68]
port 397 nsew signal input
rlabel metal2 s 357806 0 357862 800 6 la_oenb[69]
port 398 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_oenb[6]
port 399 nsew signal input
rlabel metal2 s 361118 0 361174 800 6 la_oenb[70]
port 400 nsew signal input
rlabel metal2 s 364430 0 364486 800 6 la_oenb[71]
port 401 nsew signal input
rlabel metal2 s 367742 0 367798 800 6 la_oenb[72]
port 402 nsew signal input
rlabel metal2 s 371054 0 371110 800 6 la_oenb[73]
port 403 nsew signal input
rlabel metal2 s 374366 0 374422 800 6 la_oenb[74]
port 404 nsew signal input
rlabel metal2 s 377678 0 377734 800 6 la_oenb[75]
port 405 nsew signal input
rlabel metal2 s 380990 0 381046 800 6 la_oenb[76]
port 406 nsew signal input
rlabel metal2 s 384302 0 384358 800 6 la_oenb[77]
port 407 nsew signal input
rlabel metal2 s 387614 0 387670 800 6 la_oenb[78]
port 408 nsew signal input
rlabel metal2 s 390926 0 390982 800 6 la_oenb[79]
port 409 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_oenb[7]
port 410 nsew signal input
rlabel metal2 s 394238 0 394294 800 6 la_oenb[80]
port 411 nsew signal input
rlabel metal2 s 397550 0 397606 800 6 la_oenb[81]
port 412 nsew signal input
rlabel metal2 s 400862 0 400918 800 6 la_oenb[82]
port 413 nsew signal input
rlabel metal2 s 404174 0 404230 800 6 la_oenb[83]
port 414 nsew signal input
rlabel metal2 s 407486 0 407542 800 6 la_oenb[84]
port 415 nsew signal input
rlabel metal2 s 410798 0 410854 800 6 la_oenb[85]
port 416 nsew signal input
rlabel metal2 s 414110 0 414166 800 6 la_oenb[86]
port 417 nsew signal input
rlabel metal2 s 417422 0 417478 800 6 la_oenb[87]
port 418 nsew signal input
rlabel metal2 s 420734 0 420790 800 6 la_oenb[88]
port 419 nsew signal input
rlabel metal2 s 424046 0 424102 800 6 la_oenb[89]
port 420 nsew signal input
rlabel metal2 s 155774 0 155830 800 6 la_oenb[8]
port 421 nsew signal input
rlabel metal2 s 427358 0 427414 800 6 la_oenb[90]
port 422 nsew signal input
rlabel metal2 s 430670 0 430726 800 6 la_oenb[91]
port 423 nsew signal input
rlabel metal2 s 433982 0 434038 800 6 la_oenb[92]
port 424 nsew signal input
rlabel metal2 s 437294 0 437350 800 6 la_oenb[93]
port 425 nsew signal input
rlabel metal2 s 440606 0 440662 800 6 la_oenb[94]
port 426 nsew signal input
rlabel metal2 s 443918 0 443974 800 6 la_oenb[95]
port 427 nsew signal input
rlabel metal2 s 447230 0 447286 800 6 la_oenb[96]
port 428 nsew signal input
rlabel metal2 s 450542 0 450598 800 6 la_oenb[97]
port 429 nsew signal input
rlabel metal2 s 453854 0 453910 800 6 la_oenb[98]
port 430 nsew signal input
rlabel metal2 s 457166 0 457222 800 6 la_oenb[99]
port 431 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_oenb[9]
port 432 nsew signal input
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 433 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 434 nsew ground bidirectional
rlabel metal2 s 10046 0 10102 800 6 wb_clk_i
port 435 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wb_rst_i
port 436 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_ack_o
port 437 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[0]
port 438 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 wbs_adr_i[10]
port 439 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 wbs_adr_i[11]
port 440 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_adr_i[12]
port 441 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 wbs_adr_i[13]
port 442 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_adr_i[14]
port 443 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 wbs_adr_i[15]
port 444 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_adr_i[16]
port 445 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 wbs_adr_i[17]
port 446 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 wbs_adr_i[18]
port 447 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_adr_i[19]
port 448 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[1]
port 449 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 wbs_adr_i[20]
port 450 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 wbs_adr_i[21]
port 451 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 wbs_adr_i[22]
port 452 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 wbs_adr_i[23]
port 453 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 wbs_adr_i[24]
port 454 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 wbs_adr_i[25]
port 455 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 wbs_adr_i[26]
port 456 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 wbs_adr_i[27]
port 457 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 wbs_adr_i[28]
port 458 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 wbs_adr_i[29]
port 459 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[2]
port 460 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 wbs_adr_i[30]
port 461 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 wbs_adr_i[31]
port 462 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[3]
port 463 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[4]
port 464 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[5]
port 465 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_adr_i[6]
port 466 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_adr_i[7]
port 467 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_adr_i[8]
port 468 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 wbs_adr_i[9]
port 469 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_cyc_i
port 470 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_i[0]
port 471 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 wbs_dat_i[10]
port 472 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 wbs_dat_i[11]
port 473 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_i[12]
port 474 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_i[13]
port 475 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 wbs_dat_i[14]
port 476 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_dat_i[15]
port 477 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 wbs_dat_i[16]
port 478 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 wbs_dat_i[17]
port 479 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 wbs_dat_i[18]
port 480 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 wbs_dat_i[19]
port 481 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[1]
port 482 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 wbs_dat_i[20]
port 483 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 wbs_dat_i[21]
port 484 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 wbs_dat_i[22]
port 485 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 wbs_dat_i[23]
port 486 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 wbs_dat_i[24]
port 487 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 wbs_dat_i[25]
port 488 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 wbs_dat_i[26]
port 489 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 wbs_dat_i[27]
port 490 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 wbs_dat_i[28]
port 491 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 wbs_dat_i[29]
port 492 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[2]
port 493 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 wbs_dat_i[30]
port 494 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 wbs_dat_i[31]
port 495 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[3]
port 496 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_i[4]
port 497 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_i[5]
port 498 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_dat_i[6]
port 499 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_i[7]
port 500 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_dat_i[8]
port 501 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 wbs_dat_i[9]
port 502 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[0]
port 503 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 wbs_dat_o[10]
port 504 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_o[11]
port 505 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 wbs_dat_o[12]
port 506 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 wbs_dat_o[13]
port 507 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 wbs_dat_o[14]
port 508 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 wbs_dat_o[15]
port 509 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 wbs_dat_o[16]
port 510 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_o[17]
port 511 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 wbs_dat_o[18]
port 512 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 wbs_dat_o[19]
port 513 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[1]
port 514 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 wbs_dat_o[20]
port 515 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 wbs_dat_o[21]
port 516 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 wbs_dat_o[22]
port 517 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 wbs_dat_o[23]
port 518 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 wbs_dat_o[24]
port 519 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 wbs_dat_o[25]
port 520 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 wbs_dat_o[26]
port 521 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 wbs_dat_o[27]
port 522 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 wbs_dat_o[28]
port 523 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 wbs_dat_o[29]
port 524 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_o[2]
port 525 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 wbs_dat_o[30]
port 526 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 wbs_dat_o[31]
port 527 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[3]
port 528 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_o[4]
port 529 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_o[5]
port 530 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 wbs_dat_o[6]
port 531 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 wbs_dat_o[7]
port 532 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_o[8]
port 533 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_o[9]
port 534 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_sel_i[0]
port 535 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_sel_i[1]
port 536 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_sel_i[2]
port 537 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_sel_i[3]
port 538 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_stb_i
port 539 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_we_i
port 540 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 53427234
string GDS_FILE /home/jona/Desktop/Proyecto_Final/caravan/openlane/user_analog_proj_example/runs/24_04_02_15_31/results/signoff/user_analog_proj_example.magic.gds
string GDS_START 354794
<< end >>

