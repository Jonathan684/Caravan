magic
tech sky130A
magscale 1 2
timestamp 1715159637
<< obsli1 >>
rect 13104 5159 570808 100393
<< obsm1 >>
rect 12934 8 574158 101448
<< metal2 >>
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< obsm2 >>
rect 570 536 574154 102785
rect 692 2 1650 536
rect 1874 2 2832 536
rect 3056 2 4014 536
rect 4238 2 5196 536
rect 5420 2 6378 536
rect 6602 2 7560 536
rect 7784 2 8742 536
rect 8966 2 9924 536
rect 10148 2 11106 536
rect 11330 2 12288 536
rect 12512 2 13470 536
rect 13694 2 14652 536
rect 14876 2 15834 536
rect 16058 2 17016 536
rect 17240 2 18198 536
rect 18422 2 19380 536
rect 19604 2 20562 536
rect 20786 2 21744 536
rect 21968 2 22926 536
rect 23150 2 24108 536
rect 24332 2 25290 536
rect 25514 2 26472 536
rect 26696 2 27654 536
rect 27878 2 28836 536
rect 29060 2 30018 536
rect 30242 2 31200 536
rect 31424 2 32382 536
rect 32606 2 33564 536
rect 33788 2 34746 536
rect 34970 2 35928 536
rect 36152 2 37110 536
rect 37334 2 38292 536
rect 38516 2 39474 536
rect 39698 2 40656 536
rect 40880 2 41838 536
rect 42062 2 43020 536
rect 43244 2 44202 536
rect 44426 2 45384 536
rect 45608 2 46566 536
rect 46790 2 47748 536
rect 47972 2 48930 536
rect 49154 2 50112 536
rect 50336 2 51294 536
rect 51518 2 52476 536
rect 52700 2 53658 536
rect 53882 2 54840 536
rect 55064 2 56022 536
rect 56246 2 57204 536
rect 57428 2 58386 536
rect 58610 2 59568 536
rect 59792 2 60750 536
rect 60974 2 61932 536
rect 62156 2 63114 536
rect 63338 2 64296 536
rect 64520 2 65478 536
rect 65702 2 66660 536
rect 66884 2 67842 536
rect 68066 2 69024 536
rect 69248 2 70206 536
rect 70430 2 71388 536
rect 71612 2 72570 536
rect 72794 2 73752 536
rect 73976 2 74934 536
rect 75158 2 76116 536
rect 76340 2 77298 536
rect 77522 2 78480 536
rect 78704 2 79662 536
rect 79886 2 80844 536
rect 81068 2 82026 536
rect 82250 2 83208 536
rect 83432 2 84390 536
rect 84614 2 85572 536
rect 85796 2 86754 536
rect 86978 2 87936 536
rect 88160 2 89118 536
rect 89342 2 90300 536
rect 90524 2 91482 536
rect 91706 2 92664 536
rect 92888 2 93846 536
rect 94070 2 95028 536
rect 95252 2 96210 536
rect 96434 2 97392 536
rect 97616 2 98574 536
rect 98798 2 99756 536
rect 99980 2 100938 536
rect 101162 2 102120 536
rect 102344 2 103302 536
rect 103526 2 104484 536
rect 104708 2 105666 536
rect 105890 2 106848 536
rect 107072 2 108030 536
rect 108254 2 109212 536
rect 109436 2 110394 536
rect 110618 2 111576 536
rect 111800 2 112758 536
rect 112982 2 113940 536
rect 114164 2 115122 536
rect 115346 2 116304 536
rect 116528 2 117486 536
rect 117710 2 118668 536
rect 118892 2 119850 536
rect 120074 2 121032 536
rect 121256 2 122214 536
rect 122438 2 123396 536
rect 123620 2 124578 536
rect 124802 2 125760 536
rect 125984 2 126942 536
rect 127166 2 128124 536
rect 128348 2 129306 536
rect 129530 2 130488 536
rect 130712 2 131670 536
rect 131894 2 132852 536
rect 133076 2 134034 536
rect 134258 2 135216 536
rect 135440 2 136398 536
rect 136622 2 137580 536
rect 137804 2 138762 536
rect 138986 2 139944 536
rect 140168 2 141126 536
rect 141350 2 142308 536
rect 142532 2 143490 536
rect 143714 2 144672 536
rect 144896 2 145854 536
rect 146078 2 147036 536
rect 147260 2 148218 536
rect 148442 2 149400 536
rect 149624 2 150582 536
rect 150806 2 151764 536
rect 151988 2 152946 536
rect 153170 2 154128 536
rect 154352 2 155310 536
rect 155534 2 156492 536
rect 156716 2 157674 536
rect 157898 2 158856 536
rect 159080 2 160038 536
rect 160262 2 161220 536
rect 161444 2 162402 536
rect 162626 2 163584 536
rect 163808 2 164766 536
rect 164990 2 165948 536
rect 166172 2 167130 536
rect 167354 2 168312 536
rect 168536 2 169494 536
rect 169718 2 170676 536
rect 170900 2 171858 536
rect 172082 2 173040 536
rect 173264 2 174222 536
rect 174446 2 175404 536
rect 175628 2 176586 536
rect 176810 2 177768 536
rect 177992 2 178950 536
rect 179174 2 180132 536
rect 180356 2 181314 536
rect 181538 2 182496 536
rect 182720 2 183678 536
rect 183902 2 184860 536
rect 185084 2 186042 536
rect 186266 2 187224 536
rect 187448 2 188406 536
rect 188630 2 189588 536
rect 189812 2 190770 536
rect 190994 2 191952 536
rect 192176 2 193134 536
rect 193358 2 194316 536
rect 194540 2 195498 536
rect 195722 2 196680 536
rect 196904 2 197862 536
rect 198086 2 199044 536
rect 199268 2 200226 536
rect 200450 2 201408 536
rect 201632 2 202590 536
rect 202814 2 203772 536
rect 203996 2 204954 536
rect 205178 2 206136 536
rect 206360 2 207318 536
rect 207542 2 208500 536
rect 208724 2 209682 536
rect 209906 2 210864 536
rect 211088 2 212046 536
rect 212270 2 213228 536
rect 213452 2 214410 536
rect 214634 2 215592 536
rect 215816 2 216774 536
rect 216998 2 217956 536
rect 218180 2 219138 536
rect 219362 2 220320 536
rect 220544 2 221502 536
rect 221726 2 222684 536
rect 222908 2 223866 536
rect 224090 2 225048 536
rect 225272 2 226230 536
rect 226454 2 227412 536
rect 227636 2 228594 536
rect 228818 2 229776 536
rect 230000 2 230958 536
rect 231182 2 232140 536
rect 232364 2 233322 536
rect 233546 2 234504 536
rect 234728 2 235686 536
rect 235910 2 236868 536
rect 237092 2 238050 536
rect 238274 2 239232 536
rect 239456 2 240414 536
rect 240638 2 241596 536
rect 241820 2 242778 536
rect 243002 2 243960 536
rect 244184 2 245142 536
rect 245366 2 246324 536
rect 246548 2 247506 536
rect 247730 2 248688 536
rect 248912 2 249870 536
rect 250094 2 251052 536
rect 251276 2 252234 536
rect 252458 2 253416 536
rect 253640 2 254598 536
rect 254822 2 255780 536
rect 256004 2 256962 536
rect 257186 2 258144 536
rect 258368 2 259326 536
rect 259550 2 260508 536
rect 260732 2 261690 536
rect 261914 2 262872 536
rect 263096 2 264054 536
rect 264278 2 265236 536
rect 265460 2 266418 536
rect 266642 2 267600 536
rect 267824 2 268782 536
rect 269006 2 269964 536
rect 270188 2 271146 536
rect 271370 2 272328 536
rect 272552 2 273510 536
rect 273734 2 274692 536
rect 274916 2 275874 536
rect 276098 2 277056 536
rect 277280 2 278238 536
rect 278462 2 279420 536
rect 279644 2 280602 536
rect 280826 2 281784 536
rect 282008 2 282966 536
rect 283190 2 284148 536
rect 284372 2 285330 536
rect 285554 2 286512 536
rect 286736 2 287694 536
rect 287918 2 288876 536
rect 289100 2 290058 536
rect 290282 2 291240 536
rect 291464 2 292422 536
rect 292646 2 293604 536
rect 293828 2 294786 536
rect 295010 2 295968 536
rect 296192 2 297150 536
rect 297374 2 298332 536
rect 298556 2 299514 536
rect 299738 2 300696 536
rect 300920 2 301878 536
rect 302102 2 303060 536
rect 303284 2 304242 536
rect 304466 2 305424 536
rect 305648 2 306606 536
rect 306830 2 307788 536
rect 308012 2 308970 536
rect 309194 2 310152 536
rect 310376 2 311334 536
rect 311558 2 312516 536
rect 312740 2 313698 536
rect 313922 2 314880 536
rect 315104 2 316062 536
rect 316286 2 317244 536
rect 317468 2 318426 536
rect 318650 2 319608 536
rect 319832 2 320790 536
rect 321014 2 321972 536
rect 322196 2 323154 536
rect 323378 2 324336 536
rect 324560 2 325518 536
rect 325742 2 326700 536
rect 326924 2 327882 536
rect 328106 2 329064 536
rect 329288 2 330246 536
rect 330470 2 331428 536
rect 331652 2 332610 536
rect 332834 2 333792 536
rect 334016 2 334974 536
rect 335198 2 336156 536
rect 336380 2 337338 536
rect 337562 2 338520 536
rect 338744 2 339702 536
rect 339926 2 340884 536
rect 341108 2 342066 536
rect 342290 2 343248 536
rect 343472 2 344430 536
rect 344654 2 345612 536
rect 345836 2 346794 536
rect 347018 2 347976 536
rect 348200 2 349158 536
rect 349382 2 350340 536
rect 350564 2 351522 536
rect 351746 2 352704 536
rect 352928 2 353886 536
rect 354110 2 355068 536
rect 355292 2 356250 536
rect 356474 2 357432 536
rect 357656 2 358614 536
rect 358838 2 359796 536
rect 360020 2 360978 536
rect 361202 2 362160 536
rect 362384 2 363342 536
rect 363566 2 364524 536
rect 364748 2 365706 536
rect 365930 2 366888 536
rect 367112 2 368070 536
rect 368294 2 369252 536
rect 369476 2 370434 536
rect 370658 2 371616 536
rect 371840 2 372798 536
rect 373022 2 373980 536
rect 374204 2 375162 536
rect 375386 2 376344 536
rect 376568 2 377526 536
rect 377750 2 378708 536
rect 378932 2 379890 536
rect 380114 2 381072 536
rect 381296 2 382254 536
rect 382478 2 383436 536
rect 383660 2 384618 536
rect 384842 2 385800 536
rect 386024 2 386982 536
rect 387206 2 388164 536
rect 388388 2 389346 536
rect 389570 2 390528 536
rect 390752 2 391710 536
rect 391934 2 392892 536
rect 393116 2 394074 536
rect 394298 2 395256 536
rect 395480 2 396438 536
rect 396662 2 397620 536
rect 397844 2 398802 536
rect 399026 2 399984 536
rect 400208 2 401166 536
rect 401390 2 402348 536
rect 402572 2 403530 536
rect 403754 2 404712 536
rect 404936 2 405894 536
rect 406118 2 407076 536
rect 407300 2 408258 536
rect 408482 2 409440 536
rect 409664 2 410622 536
rect 410846 2 411804 536
rect 412028 2 412986 536
rect 413210 2 414168 536
rect 414392 2 415350 536
rect 415574 2 416532 536
rect 416756 2 417714 536
rect 417938 2 418896 536
rect 419120 2 420078 536
rect 420302 2 421260 536
rect 421484 2 422442 536
rect 422666 2 423624 536
rect 423848 2 424806 536
rect 425030 2 425988 536
rect 426212 2 427170 536
rect 427394 2 428352 536
rect 428576 2 429534 536
rect 429758 2 430716 536
rect 430940 2 431898 536
rect 432122 2 433080 536
rect 433304 2 434262 536
rect 434486 2 435444 536
rect 435668 2 436626 536
rect 436850 2 437808 536
rect 438032 2 438990 536
rect 439214 2 440172 536
rect 440396 2 441354 536
rect 441578 2 442536 536
rect 442760 2 443718 536
rect 443942 2 444900 536
rect 445124 2 446082 536
rect 446306 2 447264 536
rect 447488 2 448446 536
rect 448670 2 449628 536
rect 449852 2 450810 536
rect 451034 2 451992 536
rect 452216 2 453174 536
rect 453398 2 454356 536
rect 454580 2 455538 536
rect 455762 2 456720 536
rect 456944 2 457902 536
rect 458126 2 459084 536
rect 459308 2 460266 536
rect 460490 2 461448 536
rect 461672 2 462630 536
rect 462854 2 463812 536
rect 464036 2 464994 536
rect 465218 2 466176 536
rect 466400 2 467358 536
rect 467582 2 468540 536
rect 468764 2 469722 536
rect 469946 2 470904 536
rect 471128 2 472086 536
rect 472310 2 473268 536
rect 473492 2 474450 536
rect 474674 2 475632 536
rect 475856 2 476814 536
rect 477038 2 477996 536
rect 478220 2 479178 536
rect 479402 2 480360 536
rect 480584 2 481542 536
rect 481766 2 482724 536
rect 482948 2 483906 536
rect 484130 2 485088 536
rect 485312 2 486270 536
rect 486494 2 487452 536
rect 487676 2 488634 536
rect 488858 2 489816 536
rect 490040 2 490998 536
rect 491222 2 492180 536
rect 492404 2 493362 536
rect 493586 2 494544 536
rect 494768 2 495726 536
rect 495950 2 496908 536
rect 497132 2 498090 536
rect 498314 2 499272 536
rect 499496 2 500454 536
rect 500678 2 501636 536
rect 501860 2 502818 536
rect 503042 2 504000 536
rect 504224 2 505182 536
rect 505406 2 506364 536
rect 506588 2 507546 536
rect 507770 2 508728 536
rect 508952 2 509910 536
rect 510134 2 511092 536
rect 511316 2 512274 536
rect 512498 2 513456 536
rect 513680 2 514638 536
rect 514862 2 515820 536
rect 516044 2 517002 536
rect 517226 2 518184 536
rect 518408 2 519366 536
rect 519590 2 520548 536
rect 520772 2 521730 536
rect 521954 2 522912 536
rect 523136 2 524094 536
rect 524318 2 525276 536
rect 525500 2 526458 536
rect 526682 2 527640 536
rect 527864 2 528822 536
rect 529046 2 530004 536
rect 530228 2 531186 536
rect 531410 2 532368 536
rect 532592 2 533550 536
rect 533774 2 534732 536
rect 534956 2 535914 536
rect 536138 2 537096 536
rect 537320 2 538278 536
rect 538502 2 539460 536
rect 539684 2 540642 536
rect 540866 2 541824 536
rect 542048 2 543006 536
rect 543230 2 544188 536
rect 544412 2 545370 536
rect 545594 2 546552 536
rect 546776 2 547734 536
rect 547958 2 548916 536
rect 549140 2 550098 536
rect 550322 2 551280 536
rect 551504 2 552462 536
rect 552686 2 553644 536
rect 553868 2 554826 536
rect 555050 2 556008 536
rect 556232 2 557190 536
rect 557414 2 558372 536
rect 558596 2 559554 536
rect 559778 2 560736 536
rect 560960 2 561918 536
rect 562142 2 563100 536
rect 563324 2 564282 536
rect 564506 2 565464 536
rect 565688 2 566646 536
rect 566870 2 567828 536
rect 568052 2 569010 536
rect 569234 2 570192 536
rect 570416 2 571374 536
rect 571598 2 572556 536
rect 572780 2 573738 536
rect 573962 2 574154 536
<< metal3 >>
rect 16194 702300 21194 704000
rect 68194 702300 73194 704000
rect 120194 702300 125194 704000
rect 170894 702300 173094 704000
rect 173394 702300 175594 704000
rect 175894 702300 180894 704000
rect 222594 702300 224794 704000
rect 225094 702300 227294 704000
rect 227594 702300 232594 704000
rect 324294 702300 326494 704000
rect 326794 702300 328994 704000
rect 329294 702300 334294 704000
rect 413394 702300 418394 704000
rect 465394 702300 470394 704000
rect 566594 702300 571594 704000
rect 0 680242 1700 685242
rect 582300 677984 584000 682984
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< obsm3 >>
rect 560 506722 583520 506972
rect 430 505812 583520 506722
rect 560 505540 583520 505812
rect 430 500242 583520 505540
rect 430 499970 583440 500242
rect 430 499060 583520 499970
rect 430 498788 583440 499060
rect 430 497878 583520 498788
rect 430 497606 583440 497878
rect 430 496696 583520 497606
rect 430 496424 583440 496696
rect 430 495514 583520 496424
rect 430 495242 583440 495514
rect 430 494332 583520 495242
rect 430 494060 583440 494332
rect 430 468500 583520 494060
rect 560 468228 583520 468500
rect 430 467318 583520 468228
rect 560 467046 583520 467318
rect 430 466136 583520 467046
rect 560 465864 583520 466136
rect 430 464954 583520 465864
rect 560 464682 583520 464954
rect 430 463772 583520 464682
rect 560 463500 583520 463772
rect 430 462590 583520 463500
rect 560 462318 583520 462590
rect 430 455820 583520 462318
rect 430 455548 583440 455820
rect 430 454638 583520 455548
rect 430 454366 583440 454638
rect 430 453456 583520 454366
rect 430 453184 583440 453456
rect 430 452274 583520 453184
rect 430 452002 583440 452274
rect 430 451092 583520 452002
rect 430 450820 583440 451092
rect 430 449910 583520 450820
rect 430 449638 583440 449910
rect 430 425278 583520 449638
rect 560 425006 583520 425278
rect 430 424096 583520 425006
rect 560 423824 583520 424096
rect 430 422914 583520 423824
rect 560 422642 583520 422914
rect 430 421732 583520 422642
rect 560 421460 583520 421732
rect 430 420550 583520 421460
rect 560 420278 583520 420550
rect 430 419368 583520 420278
rect 560 419096 583520 419368
rect 430 411398 583520 419096
rect 430 411126 583440 411398
rect 430 410216 583520 411126
rect 430 409944 583440 410216
rect 430 409034 583520 409944
rect 430 408762 583440 409034
rect 430 407852 583520 408762
rect 430 407580 583440 407852
rect 430 406670 583520 407580
rect 430 406398 583440 406670
rect 430 405488 583520 406398
rect 430 405216 583440 405488
rect 430 382056 583520 405216
rect 560 381784 583520 382056
rect 430 380874 583520 381784
rect 560 380602 583520 380874
rect 430 379692 583520 380602
rect 560 379420 583520 379692
rect 430 378510 583520 379420
rect 560 378238 583520 378510
rect 430 377328 583520 378238
rect 560 377056 583520 377328
rect 430 376146 583520 377056
rect 560 375874 583520 376146
rect 430 364976 583520 375874
rect 430 364704 583440 364976
rect 430 363794 583520 364704
rect 430 363522 583440 363794
rect 430 362612 583520 363522
rect 430 362340 583440 362612
rect 430 361430 583520 362340
rect 430 361158 583440 361430
rect 430 360248 583520 361158
rect 430 359976 583440 360248
rect 430 359066 583520 359976
rect 430 358794 583440 359066
rect 430 338834 583520 358794
rect 560 338562 583520 338834
rect 430 337652 583520 338562
rect 560 337380 583520 337652
rect 430 336470 583520 337380
rect 560 336198 583520 336470
rect 430 335288 583520 336198
rect 560 335016 583520 335288
rect 430 334106 583520 335016
rect 560 333834 583520 334106
rect 430 332924 583520 333834
rect 560 332652 583520 332924
rect 430 319754 583520 332652
rect 430 319482 583440 319754
rect 430 318572 583520 319482
rect 430 318300 583440 318572
rect 430 317390 583520 318300
rect 430 317118 583440 317390
rect 430 316208 583520 317118
rect 430 315936 583440 316208
rect 430 315026 583520 315936
rect 430 314754 583440 315026
rect 430 313844 583520 314754
rect 430 313572 583440 313844
rect 430 295612 583520 313572
rect 560 295340 583520 295612
rect 430 294430 583520 295340
rect 560 294158 583520 294430
rect 430 293248 583520 294158
rect 560 292976 583520 293248
rect 430 292066 583520 292976
rect 560 291794 583520 292066
rect 430 290884 583520 291794
rect 560 290612 583520 290884
rect 430 289702 583520 290612
rect 560 289430 583520 289702
rect 430 275332 583520 289430
rect 430 275060 583440 275332
rect 430 274150 583520 275060
rect 430 273878 583440 274150
rect 430 272968 583520 273878
rect 430 272696 583440 272968
rect 430 271786 583520 272696
rect 430 271514 583440 271786
rect 430 270604 583520 271514
rect 430 270332 583440 270604
rect 430 269422 583520 270332
rect 430 269150 583440 269422
rect 430 252590 583520 269150
rect 560 252318 583520 252590
rect 430 251408 583520 252318
rect 560 251136 583520 251408
rect 430 250226 583520 251136
rect 560 249954 583520 250226
rect 430 249044 583520 249954
rect 560 248772 583520 249044
rect 430 247862 583520 248772
rect 560 247590 583520 247862
rect 430 246680 583520 247590
rect 560 246408 583520 246680
rect 430 124968 583520 246408
rect 560 124696 583520 124968
rect 430 123786 583520 124696
rect 560 123514 583520 123786
rect 430 122604 583520 123514
rect 560 122332 583520 122604
rect 430 121422 583520 122332
rect 560 121150 583520 121422
rect 430 120240 583520 121150
rect 560 119968 583520 120240
rect 430 119058 583520 119968
rect 560 118786 583520 119058
rect 430 95310 583520 118786
rect 430 95038 583440 95310
rect 430 94128 583520 95038
rect 430 93856 583440 94128
rect 430 92946 583520 93856
rect 430 92674 583440 92946
rect 430 91764 583520 92674
rect 430 91492 583440 91764
rect 430 81746 583520 91492
rect 560 81474 583520 81746
rect 430 80564 583520 81474
rect 560 80292 583520 80564
rect 430 79382 583520 80292
rect 560 79110 583520 79382
rect 430 78200 583520 79110
rect 560 77928 583520 78200
rect 430 77018 583520 77928
rect 560 76746 583520 77018
rect 430 75836 583520 76746
rect 560 75564 583520 75836
rect 430 50652 583520 75564
rect 430 50380 583440 50652
rect 430 49470 583520 50380
rect 430 49198 583440 49470
rect 430 48288 583520 49198
rect 430 48016 583440 48288
rect 430 47106 583520 48016
rect 430 46834 583440 47106
rect 430 38524 583520 46834
rect 560 38252 583520 38524
rect 430 37342 583520 38252
rect 560 37070 583520 37342
rect 430 36160 583520 37070
rect 560 35888 583520 36160
rect 430 34978 583520 35888
rect 560 34706 583520 34978
rect 430 33796 583520 34706
rect 560 33524 583520 33796
rect 430 32614 583520 33524
rect 560 32342 583520 32614
rect 430 24194 583520 32342
rect 430 23922 583440 24194
rect 430 23012 583520 23922
rect 430 22740 583440 23012
rect 430 21830 583520 22740
rect 430 21558 583440 21830
rect 430 20648 583520 21558
rect 430 20376 583440 20648
rect 430 19466 583520 20376
rect 430 19194 583440 19466
rect 430 18284 583520 19194
rect 430 18012 583440 18284
rect 430 17102 583520 18012
rect 560 16830 583440 17102
rect 430 15920 583520 16830
rect 560 15648 583440 15920
rect 430 14738 583520 15648
rect 560 14466 583440 14738
rect 430 13556 583520 14466
rect 560 13284 583440 13556
rect 430 12374 583520 13284
rect 560 12102 583440 12374
rect 430 11192 583520 12102
rect 560 10920 583440 11192
rect 430 10010 583520 10920
rect 560 9738 583440 10010
rect 430 8828 583520 9738
rect 560 8556 583440 8828
rect 430 7646 583520 8556
rect 560 7374 583440 7646
rect 430 6464 583520 7374
rect 560 6192 583440 6464
rect 430 5282 583520 6192
rect 560 5010 583440 5282
rect 430 4100 583520 5010
rect 560 3828 583440 4100
rect 430 2918 583520 3828
rect 560 2646 583440 2918
rect 430 1736 583520 2646
rect 560 1464 583440 1736
rect 430 35 583520 1464
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -7654 2414 711590
rect 5514 -7654 6134 711590
rect 9234 -7654 9854 711590
rect 12954 -7654 13574 711590
rect 16674 -7654 17294 711590
rect 20394 -7654 21014 711590
rect 24114 -7654 24734 711590
rect 27834 -7654 28454 711590
rect 37794 -7654 38414 711590
rect 41514 -7654 42134 711590
rect 45234 -7654 45854 711590
rect 48954 -7654 49574 711590
rect 52674 -7654 53294 711590
rect 56394 -7654 57014 711590
rect 60114 -7654 60734 711590
rect 63834 -7654 64454 711590
rect 73794 -7654 74414 711590
rect 77514 102564 78134 711590
rect 81234 -7654 81854 711590
rect 84954 -7654 85574 711590
rect 88674 -7654 89294 711590
rect 92394 102564 93014 711590
rect 96114 -7654 96734 711590
rect 99834 -7654 100454 711590
rect 109794 -7654 110414 711590
rect 113514 -7654 114134 711590
rect 117234 -7654 117854 711590
rect 120954 -7654 121574 711590
rect 124674 -7654 125294 711590
rect 128394 -7654 129014 711590
rect 132114 -7654 132734 711590
rect 135834 -7654 136454 711590
rect 145794 -7654 146414 711590
rect 149514 -7654 150134 711590
rect 153234 -7654 153854 711590
rect 156954 -7654 157574 711590
rect 160674 -7654 161294 711590
rect 164394 -7654 165014 711590
rect 168114 -7654 168734 711590
rect 171834 -7654 172454 711590
rect 181794 -7654 182414 711590
rect 185514 102564 186134 711590
rect 189234 -7654 189854 711590
rect 192954 -7654 193574 711590
rect 196674 -7654 197294 711590
rect 200394 102564 201014 711590
rect 204114 -7654 204734 711590
rect 207834 -7654 208454 711590
rect 217794 -7654 218414 711590
rect 221514 -7654 222134 711590
rect 225234 -7654 225854 711590
rect 228954 -7654 229574 711590
rect 232674 -7654 233294 711590
rect 236394 -7654 237014 711590
rect 240114 -7654 240734 711590
rect 243834 -7654 244454 711590
rect 253794 -7654 254414 711590
rect 257514 -7654 258134 711590
rect 261234 102564 261854 711590
rect 264954 -7654 265574 711590
rect 268674 -7654 269294 711590
rect 272394 -7654 273014 711590
rect 276114 -7654 276734 711590
rect 279834 -7654 280454 711590
rect 289794 -7654 290414 711590
rect 293514 -7654 294134 711590
rect 297234 -7654 297854 711590
rect 300954 -7654 301574 711590
rect 304674 -7654 305294 711590
rect 308394 102564 309014 711590
rect 312114 -7654 312734 711590
rect 315834 -7654 316454 711590
rect 325794 -7654 326414 711590
rect 329514 -7654 330134 711590
rect 333234 -7654 333854 711590
rect 336954 -7654 337574 711590
rect 340674 -7654 341294 711590
rect 344394 -7654 345014 711590
rect 348114 -7654 348734 711590
rect 351834 -7654 352454 711590
rect 361794 -7654 362414 711590
rect 365514 -7654 366134 711590
rect 369234 102564 369854 711590
rect 372954 -7654 373574 711590
rect 376674 -7654 377294 711590
rect 380394 -7654 381014 711590
rect 384114 102564 384734 711590
rect 387834 -7654 388454 711590
rect 397794 -7654 398414 711590
rect 401514 -7654 402134 711590
rect 405234 -7654 405854 711590
rect 408954 -7654 409574 711590
rect 412674 -7654 413294 711590
rect 416394 -7654 417014 711590
rect 420114 -7654 420734 711590
rect 423834 -7654 424454 711590
rect 433794 -7654 434414 711590
rect 437514 -7654 438134 711590
rect 441234 -7654 441854 711590
rect 444954 -7654 445574 711590
rect 448674 -7654 449294 711590
rect 452394 -7654 453014 711590
rect 456114 -7654 456734 711590
rect 459834 -7654 460454 711590
rect 469794 -7654 470414 711590
rect 473514 -7654 474134 711590
rect 477234 102564 477854 711590
rect 480954 -7654 481574 711590
rect 484674 -7654 485294 711590
rect 488394 -7654 489014 711590
rect 492114 102564 492734 711590
rect 495834 -7654 496454 711590
rect 505794 -7654 506414 711590
rect 509514 -7654 510134 711590
rect 513234 -7654 513854 711590
rect 516954 -7654 517574 711590
rect 520674 -7654 521294 711590
rect 524394 -7654 525014 711590
rect 528114 -7654 528734 711590
rect 531834 -7654 532454 711590
rect 541794 -7654 542414 711590
rect 545514 -7654 546134 711590
rect 549234 -7654 549854 711590
rect 552954 -7654 553574 711590
rect 556674 -7654 557294 711590
rect 560394 -7654 561014 711590
rect 564114 -7654 564734 711590
rect 567834 -7654 568454 711590
rect 577794 -7654 578414 711590
rect 581514 -7654 582134 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 3371 443 5434 506973
rect 6214 443 9154 506973
rect 9934 443 12874 506973
rect 13654 443 16594 506973
rect 17374 443 20314 506973
rect 21094 443 24034 506973
rect 24814 443 27754 506973
rect 28534 443 37714 506973
rect 38494 443 41434 506973
rect 42214 443 45154 506973
rect 45934 443 48874 506973
rect 49654 443 52594 506973
rect 53374 443 56314 506973
rect 57094 443 60034 506973
rect 60814 443 63754 506973
rect 64534 443 73714 506973
rect 74494 102484 77434 506973
rect 78214 102484 81154 506973
rect 74494 443 81154 102484
rect 81934 443 84874 506973
rect 85654 443 88594 506973
rect 89374 102484 92314 506973
rect 93094 102484 96034 506973
rect 89374 443 96034 102484
rect 96814 443 99754 506973
rect 100534 443 109714 506973
rect 110494 443 113434 506973
rect 114214 443 117154 506973
rect 117934 443 120874 506973
rect 121654 443 124594 506973
rect 125374 443 128314 506973
rect 129094 443 132034 506973
rect 132814 443 135754 506973
rect 136534 443 145714 506973
rect 146494 443 149434 506973
rect 150214 443 153154 506973
rect 153934 443 156874 506973
rect 157654 443 160594 506973
rect 161374 443 164314 506973
rect 165094 443 168034 506973
rect 168814 443 171754 506973
rect 172534 443 181714 506973
rect 182494 102484 185434 506973
rect 186214 102484 189154 506973
rect 182494 443 189154 102484
rect 189934 443 192874 506973
rect 193654 443 196594 506973
rect 197374 102484 200314 506973
rect 201094 102484 204034 506973
rect 197374 443 204034 102484
rect 204814 443 207754 506973
rect 208534 443 217714 506973
rect 218494 443 221434 506973
rect 222214 443 225154 506973
rect 225934 443 228874 506973
rect 229654 443 232594 506973
rect 233374 443 236314 506973
rect 237094 443 240034 506973
rect 240814 443 243754 506973
rect 244534 443 253714 506973
rect 254494 443 257434 506973
rect 258214 102484 261154 506973
rect 261934 102484 264874 506973
rect 258214 443 264874 102484
rect 265654 443 268594 506973
rect 269374 443 272314 506973
rect 273094 443 276034 506973
rect 276814 443 279754 506973
rect 280534 443 289714 506973
rect 290494 443 293434 506973
rect 294214 443 297154 506973
rect 297934 443 300874 506973
rect 301654 443 304594 506973
rect 305374 102484 308314 506973
rect 309094 102484 312034 506973
rect 305374 443 312034 102484
rect 312814 443 315754 506973
rect 316534 443 325714 506973
rect 326494 443 329434 506973
rect 330214 443 333154 506973
rect 333934 443 336874 506973
rect 337654 443 340594 506973
rect 341374 443 344314 506973
rect 345094 443 348034 506973
rect 348814 443 351754 506973
rect 352534 443 361714 506973
rect 362494 443 365434 506973
rect 366214 102484 369154 506973
rect 369934 102484 372874 506973
rect 366214 443 372874 102484
rect 373654 443 376594 506973
rect 377374 443 380314 506973
rect 381094 102484 384034 506973
rect 384814 102484 387754 506973
rect 381094 443 387754 102484
rect 388534 443 397714 506973
rect 398494 443 401434 506973
rect 402214 443 405154 506973
rect 405934 443 408874 506973
rect 409654 443 412594 506973
rect 413374 443 416314 506973
rect 417094 443 420034 506973
rect 420814 443 423754 506973
rect 424534 443 433714 506973
rect 434494 443 437434 506973
rect 438214 443 441154 506973
rect 441934 443 444874 506973
rect 445654 443 448594 506973
rect 449374 443 452314 506973
rect 453094 443 456034 506973
rect 456814 443 459754 506973
rect 460534 443 469714 506973
rect 470494 443 473434 506973
rect 474214 102484 477154 506973
rect 477934 102484 480874 506973
rect 474214 443 480874 102484
rect 481654 443 484594 506973
rect 485374 443 488314 506973
rect 489094 102484 492034 506973
rect 492814 102484 495754 506973
rect 489094 443 495754 102484
rect 496534 443 505714 506973
rect 506494 443 509434 506973
rect 510214 443 513154 506973
rect 513934 443 516874 506973
rect 517654 443 520594 506973
rect 521374 443 524314 506973
rect 525094 443 528034 506973
rect 528814 443 531754 506973
rect 532534 443 541714 506973
rect 542494 443 545434 506973
rect 546214 443 549154 506973
rect 549934 443 552874 506973
rect 553654 443 556594 506973
rect 557374 443 560314 506973
rect 561094 443 564034 506973
rect 564814 443 567754 506973
rect 568534 443 577714 506973
rect 578494 443 580277 506973
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -8726 694306 592650 694926
rect -8726 690586 592650 691206
rect -8726 686866 592650 687486
rect -8726 676906 592650 677526
rect -8726 673186 592650 673806
rect -8726 669466 592650 670086
rect -8726 665746 592650 666366
rect -8726 662026 592650 662646
rect -8726 658306 592650 658926
rect -8726 654586 592650 655206
rect -8726 650866 592650 651486
rect -8726 640906 592650 641526
rect -8726 637186 592650 637806
rect -8726 633466 592650 634086
rect -8726 629746 592650 630366
rect -8726 626026 592650 626646
rect -8726 622306 592650 622926
rect -8726 618586 592650 619206
rect -8726 614866 592650 615486
rect -8726 604906 592650 605526
rect -8726 601186 592650 601806
rect -8726 597466 592650 598086
rect -8726 593746 592650 594366
rect -8726 590026 592650 590646
rect -8726 586306 592650 586926
rect -8726 582586 592650 583206
rect -8726 578866 592650 579486
rect -8726 568906 592650 569526
rect -8726 565186 592650 565806
rect -8726 561466 592650 562086
rect -8726 557746 592650 558366
rect -8726 554026 592650 554646
rect -8726 550306 592650 550926
rect -8726 546586 592650 547206
rect -8726 542866 592650 543486
rect -8726 532906 592650 533526
rect -8726 529186 592650 529806
rect -8726 525466 592650 526086
rect -8726 521746 592650 522366
rect -8726 518026 592650 518646
rect -8726 514306 592650 514926
rect -8726 510586 592650 511206
rect -8726 506866 592650 507486
rect -8726 496906 592650 497526
rect -8726 493186 592650 493806
rect -8726 489466 592650 490086
rect -8726 485746 592650 486366
rect -8726 482026 592650 482646
rect -8726 478306 592650 478926
rect -8726 474586 592650 475206
rect -8726 470866 592650 471486
rect -8726 460906 592650 461526
rect -8726 457186 592650 457806
rect -8726 453466 592650 454086
rect -8726 449746 592650 450366
rect -8726 446026 592650 446646
rect -8726 442306 592650 442926
rect -8726 438586 592650 439206
rect -8726 434866 592650 435486
rect -8726 424906 592650 425526
rect -8726 421186 592650 421806
rect -8726 417466 592650 418086
rect -8726 413746 592650 414366
rect -8726 410026 592650 410646
rect -8726 406306 592650 406926
rect -8726 402586 592650 403206
rect -8726 398866 592650 399486
rect -8726 388906 592650 389526
rect -8726 385186 592650 385806
rect -8726 381466 592650 382086
rect -8726 377746 592650 378366
rect -8726 374026 592650 374646
rect -8726 370306 592650 370926
rect -8726 366586 592650 367206
rect -8726 362866 592650 363486
rect -8726 352906 592650 353526
rect -8726 349186 592650 349806
rect -8726 345466 592650 346086
rect -8726 341746 592650 342366
rect -8726 338026 592650 338646
rect -8726 334306 592650 334926
rect -8726 330586 592650 331206
rect -8726 326866 592650 327486
rect -8726 316906 592650 317526
rect -8726 313186 592650 313806
rect -8726 309466 592650 310086
rect -8726 305746 592650 306366
rect -8726 302026 592650 302646
rect -8726 298306 592650 298926
rect -8726 294586 592650 295206
rect -8726 290866 592650 291486
rect -8726 280906 592650 281526
rect -8726 277186 592650 277806
rect -8726 273466 592650 274086
rect -8726 269746 592650 270366
rect -8726 266026 592650 266646
rect -8726 262306 592650 262926
rect -8726 258586 592650 259206
rect -8726 254866 592650 255486
rect -8726 244906 592650 245526
rect -8726 241186 592650 241806
rect -8726 237466 592650 238086
rect -8726 233746 592650 234366
rect -8726 230026 592650 230646
rect -8726 226306 592650 226926
rect -8726 222586 592650 223206
rect -8726 218866 592650 219486
rect -8726 208906 592650 209526
rect -8726 205186 592650 205806
rect -8726 201466 592650 202086
rect -8726 197746 592650 198366
rect -8726 194026 592650 194646
rect -8726 190306 592650 190926
rect -8726 186586 592650 187206
rect -8726 182866 592650 183486
rect -8726 172906 592650 173526
rect -8726 169186 592650 169806
rect -8726 165466 592650 166086
rect -8726 161746 592650 162366
rect -8726 158026 592650 158646
rect -8726 154306 592650 154926
rect -8726 150586 592650 151206
rect -8726 146866 592650 147486
rect -8726 136906 592650 137526
rect -8726 133186 592650 133806
rect -8726 129466 592650 130086
rect -8726 125746 592650 126366
rect -8726 122026 592650 122646
rect -8726 118306 592650 118926
rect -8726 114586 592650 115206
rect -8726 110866 592650 111486
rect -8726 100906 592650 101526
rect -8726 97186 592650 97806
rect -8726 93466 592650 94086
rect -8726 89746 592650 90366
rect -8726 86026 592650 86646
rect -8726 82306 592650 82926
rect -8726 78586 592650 79206
rect -8726 74866 592650 75486
rect -8726 64906 592650 65526
rect -8726 61186 592650 61806
rect -8726 57466 592650 58086
rect -8726 53746 592650 54366
rect -8726 50026 592650 50646
rect -8726 46306 592650 46926
rect -8726 42586 592650 43206
rect -8726 38866 592650 39486
rect -8726 28906 592650 29526
rect -8726 25186 592650 25806
rect -8726 21466 592650 22086
rect -8726 17746 592650 18366
rect -8726 14026 592650 14646
rect -8726 10306 592650 10926
rect -8726 6586 592650 7206
rect -8726 2866 592650 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 269230 584800 269342 6 gpio_analog[0]
port 1 nsew signal bidirectional
rlabel metal3 s -800 381864 480 381976 4 gpio_analog[10]
port 2 nsew signal bidirectional
rlabel metal3 s -800 338642 480 338754 4 gpio_analog[11]
port 3 nsew signal bidirectional
rlabel metal3 s -800 295420 480 295532 4 gpio_analog[12]
port 4 nsew signal bidirectional
rlabel metal3 s -800 252398 480 252510 4 gpio_analog[13]
port 5 nsew signal bidirectional
rlabel metal3 s -800 124776 480 124888 4 gpio_analog[14]
port 6 nsew signal bidirectional
rlabel metal3 s -800 81554 480 81666 4 gpio_analog[15]
port 7 nsew signal bidirectional
rlabel metal3 s -800 38332 480 38444 4 gpio_analog[16]
port 8 nsew signal bidirectional
rlabel metal3 s -800 16910 480 17022 4 gpio_analog[17]
port 9 nsew signal bidirectional
rlabel metal3 s 583520 313652 584800 313764 6 gpio_analog[1]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 358874 584800 358986 6 gpio_analog[2]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 405296 584800 405408 6 gpio_analog[3]
port 12 nsew signal bidirectional
rlabel metal3 s 583520 449718 584800 449830 6 gpio_analog[4]
port 13 nsew signal bidirectional
rlabel metal3 s 583520 494140 584800 494252 6 gpio_analog[5]
port 14 nsew signal bidirectional
rlabel metal3 s 583520 583562 584800 583674 6 gpio_analog[6]
port 15 nsew signal bidirectional
rlabel metal3 s -800 511530 480 511642 4 gpio_analog[7]
port 16 nsew signal bidirectional
rlabel metal3 s -800 468308 480 468420 4 gpio_analog[8]
port 17 nsew signal bidirectional
rlabel metal3 s -800 425086 480 425198 4 gpio_analog[9]
port 18 nsew signal bidirectional
rlabel metal3 s 583520 270412 584800 270524 6 gpio_noesd[0]
port 19 nsew signal bidirectional
rlabel metal3 s -800 380682 480 380794 4 gpio_noesd[10]
port 20 nsew signal bidirectional
rlabel metal3 s -800 337460 480 337572 4 gpio_noesd[11]
port 21 nsew signal bidirectional
rlabel metal3 s -800 294238 480 294350 4 gpio_noesd[12]
port 22 nsew signal bidirectional
rlabel metal3 s -800 251216 480 251328 4 gpio_noesd[13]
port 23 nsew signal bidirectional
rlabel metal3 s -800 123594 480 123706 4 gpio_noesd[14]
port 24 nsew signal bidirectional
rlabel metal3 s -800 80372 480 80484 4 gpio_noesd[15]
port 25 nsew signal bidirectional
rlabel metal3 s -800 37150 480 37262 4 gpio_noesd[16]
port 26 nsew signal bidirectional
rlabel metal3 s -800 15728 480 15840 4 gpio_noesd[17]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 314834 584800 314946 6 gpio_noesd[1]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 360056 584800 360168 6 gpio_noesd[2]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 406478 584800 406590 6 gpio_noesd[3]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 450900 584800 451012 6 gpio_noesd[4]
port 31 nsew signal bidirectional
rlabel metal3 s 583520 495322 584800 495434 6 gpio_noesd[5]
port 32 nsew signal bidirectional
rlabel metal3 s 583520 584744 584800 584856 6 gpio_noesd[6]
port 33 nsew signal bidirectional
rlabel metal3 s -800 510348 480 510460 4 gpio_noesd[7]
port 34 nsew signal bidirectional
rlabel metal3 s -800 467126 480 467238 4 gpio_noesd[8]
port 35 nsew signal bidirectional
rlabel metal3 s -800 423904 480 424016 4 gpio_noesd[9]
port 36 nsew signal bidirectional
rlabel metal3 s 582300 677984 584000 682984 6 io_analog[0]
port 37 nsew signal bidirectional
rlabel metal3 s 0 680242 1700 685242 6 io_analog[10]
port 38 nsew signal bidirectional
rlabel metal3 s 566594 702300 571594 704000 6 io_analog[1]
port 39 nsew signal bidirectional
rlabel metal3 s 465394 702300 470394 704000 6 io_analog[2]
port 40 nsew signal bidirectional
rlabel metal3 s 413394 702300 418394 704000 6 io_analog[3]
port 41 nsew signal bidirectional
rlabel metal3 s 329294 702300 334294 704000 6 io_analog[4]
port 42 nsew signal bidirectional
rlabel metal3 s 227594 702300 232594 704000 6 io_analog[5]
port 43 nsew signal bidirectional
rlabel metal3 s 175894 702300 180894 704000 6 io_analog[6]
port 44 nsew signal bidirectional
rlabel metal3 s 120194 702300 125194 704000 6 io_analog[7]
port 45 nsew signal bidirectional
rlabel metal3 s 68194 702300 73194 704000 6 io_analog[8]
port 46 nsew signal bidirectional
rlabel metal3 s 16194 702300 21194 704000 6 io_analog[9]
port 47 nsew signal bidirectional
rlabel metal3 s 326794 702300 328994 704000 6 io_clamp_high[0]
port 48 nsew signal bidirectional
rlabel metal3 s 225094 702300 227294 704000 6 io_clamp_high[1]
port 49 nsew signal bidirectional
rlabel metal3 s 173394 702300 175594 704000 6 io_clamp_high[2]
port 50 nsew signal bidirectional
rlabel metal3 s 324294 702300 326494 704000 6 io_clamp_low[0]
port 51 nsew signal bidirectional
rlabel metal3 s 222594 702300 224794 704000 6 io_clamp_low[1]
port 52 nsew signal bidirectional
rlabel metal3 s 170894 702300 173094 704000 6 io_clamp_low[2]
port 53 nsew signal bidirectional
rlabel metal3 s 583520 2726 584800 2838 6 io_in[0]
port 54 nsew signal input
rlabel metal3 s 583520 408842 584800 408954 6 io_in[10]
port 55 nsew signal input
rlabel metal3 s 583520 453264 584800 453376 6 io_in[11]
port 56 nsew signal input
rlabel metal3 s 583520 497686 584800 497798 6 io_in[12]
port 57 nsew signal input
rlabel metal3 s 583520 587108 584800 587220 6 io_in[13]
port 58 nsew signal input
rlabel metal3 s -800 507984 480 508096 4 io_in[14]
port 59 nsew signal input
rlabel metal3 s -800 464762 480 464874 4 io_in[15]
port 60 nsew signal input
rlabel metal3 s -800 421540 480 421652 4 io_in[16]
port 61 nsew signal input
rlabel metal3 s -800 378318 480 378430 4 io_in[17]
port 62 nsew signal input
rlabel metal3 s -800 335096 480 335208 4 io_in[18]
port 63 nsew signal input
rlabel metal3 s -800 291874 480 291986 4 io_in[19]
port 64 nsew signal input
rlabel metal3 s 583520 7454 584800 7566 6 io_in[1]
port 65 nsew signal input
rlabel metal3 s -800 248852 480 248964 4 io_in[20]
port 66 nsew signal input
rlabel metal3 s -800 121230 480 121342 4 io_in[21]
port 67 nsew signal input
rlabel metal3 s -800 78008 480 78120 4 io_in[22]
port 68 nsew signal input
rlabel metal3 s -800 34786 480 34898 4 io_in[23]
port 69 nsew signal input
rlabel metal3 s -800 13364 480 13476 4 io_in[24]
port 70 nsew signal input
rlabel metal3 s -800 8636 480 8748 4 io_in[25]
port 71 nsew signal input
rlabel metal3 s -800 3908 480 4020 4 io_in[26]
port 72 nsew signal input
rlabel metal3 s 583520 12182 584800 12294 6 io_in[2]
port 73 nsew signal input
rlabel metal3 s 583520 16910 584800 17022 6 io_in[3]
port 74 nsew signal input
rlabel metal3 s 583520 21638 584800 21750 6 io_in[4]
port 75 nsew signal input
rlabel metal3 s 583520 48096 584800 48208 6 io_in[5]
port 76 nsew signal input
rlabel metal3 s 583520 92754 584800 92866 6 io_in[6]
port 77 nsew signal input
rlabel metal3 s 583520 272776 584800 272888 6 io_in[7]
port 78 nsew signal input
rlabel metal3 s 583520 317198 584800 317310 6 io_in[8]
port 79 nsew signal input
rlabel metal3 s 583520 362420 584800 362532 6 io_in[9]
port 80 nsew signal input
rlabel metal3 s 583520 1544 584800 1656 6 io_in_3v3[0]
port 81 nsew signal input
rlabel metal3 s 583520 407660 584800 407772 6 io_in_3v3[10]
port 82 nsew signal input
rlabel metal3 s 583520 452082 584800 452194 6 io_in_3v3[11]
port 83 nsew signal input
rlabel metal3 s 583520 496504 584800 496616 6 io_in_3v3[12]
port 84 nsew signal input
rlabel metal3 s 583520 585926 584800 586038 6 io_in_3v3[13]
port 85 nsew signal input
rlabel metal3 s -800 509166 480 509278 4 io_in_3v3[14]
port 86 nsew signal input
rlabel metal3 s -800 465944 480 466056 4 io_in_3v3[15]
port 87 nsew signal input
rlabel metal3 s -800 422722 480 422834 4 io_in_3v3[16]
port 88 nsew signal input
rlabel metal3 s -800 379500 480 379612 4 io_in_3v3[17]
port 89 nsew signal input
rlabel metal3 s -800 336278 480 336390 4 io_in_3v3[18]
port 90 nsew signal input
rlabel metal3 s -800 293056 480 293168 4 io_in_3v3[19]
port 91 nsew signal input
rlabel metal3 s 583520 6272 584800 6384 6 io_in_3v3[1]
port 92 nsew signal input
rlabel metal3 s -800 250034 480 250146 4 io_in_3v3[20]
port 93 nsew signal input
rlabel metal3 s -800 122412 480 122524 4 io_in_3v3[21]
port 94 nsew signal input
rlabel metal3 s -800 79190 480 79302 4 io_in_3v3[22]
port 95 nsew signal input
rlabel metal3 s -800 35968 480 36080 4 io_in_3v3[23]
port 96 nsew signal input
rlabel metal3 s -800 14546 480 14658 4 io_in_3v3[24]
port 97 nsew signal input
rlabel metal3 s -800 9818 480 9930 4 io_in_3v3[25]
port 98 nsew signal input
rlabel metal3 s -800 5090 480 5202 4 io_in_3v3[26]
port 99 nsew signal input
rlabel metal3 s 583520 11000 584800 11112 6 io_in_3v3[2]
port 100 nsew signal input
rlabel metal3 s 583520 15728 584800 15840 6 io_in_3v3[3]
port 101 nsew signal input
rlabel metal3 s 583520 20456 584800 20568 6 io_in_3v3[4]
port 102 nsew signal input
rlabel metal3 s 583520 46914 584800 47026 6 io_in_3v3[5]
port 103 nsew signal input
rlabel metal3 s 583520 91572 584800 91684 6 io_in_3v3[6]
port 104 nsew signal input
rlabel metal3 s 583520 271594 584800 271706 6 io_in_3v3[7]
port 105 nsew signal input
rlabel metal3 s 583520 316016 584800 316128 6 io_in_3v3[8]
port 106 nsew signal input
rlabel metal3 s 583520 361238 584800 361350 6 io_in_3v3[9]
port 107 nsew signal input
rlabel metal3 s 583520 5090 584800 5202 6 io_oeb[0]
port 108 nsew signal output
rlabel metal3 s 583520 411206 584800 411318 6 io_oeb[10]
port 109 nsew signal output
rlabel metal3 s 583520 455628 584800 455740 6 io_oeb[11]
port 110 nsew signal output
rlabel metal3 s 583520 500050 584800 500162 6 io_oeb[12]
port 111 nsew signal output
rlabel metal3 s 583520 589472 584800 589584 6 io_oeb[13]
port 112 nsew signal output
rlabel metal3 s -800 505620 480 505732 4 io_oeb[14]
port 113 nsew signal output
rlabel metal3 s -800 462398 480 462510 4 io_oeb[15]
port 114 nsew signal output
rlabel metal3 s -800 419176 480 419288 4 io_oeb[16]
port 115 nsew signal output
rlabel metal3 s -800 375954 480 376066 4 io_oeb[17]
port 116 nsew signal output
rlabel metal3 s -800 332732 480 332844 4 io_oeb[18]
port 117 nsew signal output
rlabel metal3 s -800 289510 480 289622 4 io_oeb[19]
port 118 nsew signal output
rlabel metal3 s 583520 9818 584800 9930 6 io_oeb[1]
port 119 nsew signal output
rlabel metal3 s -800 246488 480 246600 4 io_oeb[20]
port 120 nsew signal output
rlabel metal3 s -800 118866 480 118978 4 io_oeb[21]
port 121 nsew signal output
rlabel metal3 s -800 75644 480 75756 4 io_oeb[22]
port 122 nsew signal output
rlabel metal3 s -800 32422 480 32534 4 io_oeb[23]
port 123 nsew signal output
rlabel metal3 s -800 11000 480 11112 4 io_oeb[24]
port 124 nsew signal output
rlabel metal3 s -800 6272 480 6384 4 io_oeb[25]
port 125 nsew signal output
rlabel metal3 s -800 1544 480 1656 4 io_oeb[26]
port 126 nsew signal output
rlabel metal3 s 583520 14546 584800 14658 6 io_oeb[2]
port 127 nsew signal output
rlabel metal3 s 583520 19274 584800 19386 6 io_oeb[3]
port 128 nsew signal output
rlabel metal3 s 583520 24002 584800 24114 6 io_oeb[4]
port 129 nsew signal output
rlabel metal3 s 583520 50460 584800 50572 6 io_oeb[5]
port 130 nsew signal output
rlabel metal3 s 583520 95118 584800 95230 6 io_oeb[6]
port 131 nsew signal output
rlabel metal3 s 583520 275140 584800 275252 6 io_oeb[7]
port 132 nsew signal output
rlabel metal3 s 583520 319562 584800 319674 6 io_oeb[8]
port 133 nsew signal output
rlabel metal3 s 583520 364784 584800 364896 6 io_oeb[9]
port 134 nsew signal output
rlabel metal3 s 583520 3908 584800 4020 6 io_out[0]
port 135 nsew signal output
rlabel metal3 s 583520 410024 584800 410136 6 io_out[10]
port 136 nsew signal output
rlabel metal3 s 583520 454446 584800 454558 6 io_out[11]
port 137 nsew signal output
rlabel metal3 s 583520 498868 584800 498980 6 io_out[12]
port 138 nsew signal output
rlabel metal3 s 583520 588290 584800 588402 6 io_out[13]
port 139 nsew signal output
rlabel metal3 s -800 506802 480 506914 4 io_out[14]
port 140 nsew signal output
rlabel metal3 s -800 463580 480 463692 4 io_out[15]
port 141 nsew signal output
rlabel metal3 s -800 420358 480 420470 4 io_out[16]
port 142 nsew signal output
rlabel metal3 s -800 377136 480 377248 4 io_out[17]
port 143 nsew signal output
rlabel metal3 s -800 333914 480 334026 4 io_out[18]
port 144 nsew signal output
rlabel metal3 s -800 290692 480 290804 4 io_out[19]
port 145 nsew signal output
rlabel metal3 s 583520 8636 584800 8748 6 io_out[1]
port 146 nsew signal output
rlabel metal3 s -800 247670 480 247782 4 io_out[20]
port 147 nsew signal output
rlabel metal3 s -800 120048 480 120160 4 io_out[21]
port 148 nsew signal output
rlabel metal3 s -800 76826 480 76938 4 io_out[22]
port 149 nsew signal output
rlabel metal3 s -800 33604 480 33716 4 io_out[23]
port 150 nsew signal output
rlabel metal3 s -800 12182 480 12294 4 io_out[24]
port 151 nsew signal output
rlabel metal3 s -800 7454 480 7566 4 io_out[25]
port 152 nsew signal output
rlabel metal3 s -800 2726 480 2838 4 io_out[26]
port 153 nsew signal output
rlabel metal3 s 583520 13364 584800 13476 6 io_out[2]
port 154 nsew signal output
rlabel metal3 s 583520 18092 584800 18204 6 io_out[3]
port 155 nsew signal output
rlabel metal3 s 583520 22820 584800 22932 6 io_out[4]
port 156 nsew signal output
rlabel metal3 s 583520 49278 584800 49390 6 io_out[5]
port 157 nsew signal output
rlabel metal3 s 583520 93936 584800 94048 6 io_out[6]
port 158 nsew signal output
rlabel metal3 s 583520 273958 584800 274070 6 io_out[7]
port 159 nsew signal output
rlabel metal3 s 583520 318380 584800 318492 6 io_out[8]
port 160 nsew signal output
rlabel metal3 s 583520 363602 584800 363714 6 io_out[9]
port 161 nsew signal output
rlabel metal2 s 125816 -800 125928 480 8 la_data_in[0]
port 162 nsew signal input
rlabel metal2 s 480416 -800 480528 480 8 la_data_in[100]
port 163 nsew signal input
rlabel metal2 s 483962 -800 484074 480 8 la_data_in[101]
port 164 nsew signal input
rlabel metal2 s 487508 -800 487620 480 8 la_data_in[102]
port 165 nsew signal input
rlabel metal2 s 491054 -800 491166 480 8 la_data_in[103]
port 166 nsew signal input
rlabel metal2 s 494600 -800 494712 480 8 la_data_in[104]
port 167 nsew signal input
rlabel metal2 s 498146 -800 498258 480 8 la_data_in[105]
port 168 nsew signal input
rlabel metal2 s 501692 -800 501804 480 8 la_data_in[106]
port 169 nsew signal input
rlabel metal2 s 505238 -800 505350 480 8 la_data_in[107]
port 170 nsew signal input
rlabel metal2 s 508784 -800 508896 480 8 la_data_in[108]
port 171 nsew signal input
rlabel metal2 s 512330 -800 512442 480 8 la_data_in[109]
port 172 nsew signal input
rlabel metal2 s 161276 -800 161388 480 8 la_data_in[10]
port 173 nsew signal input
rlabel metal2 s 515876 -800 515988 480 8 la_data_in[110]
port 174 nsew signal input
rlabel metal2 s 519422 -800 519534 480 8 la_data_in[111]
port 175 nsew signal input
rlabel metal2 s 522968 -800 523080 480 8 la_data_in[112]
port 176 nsew signal input
rlabel metal2 s 526514 -800 526626 480 8 la_data_in[113]
port 177 nsew signal input
rlabel metal2 s 530060 -800 530172 480 8 la_data_in[114]
port 178 nsew signal input
rlabel metal2 s 533606 -800 533718 480 8 la_data_in[115]
port 179 nsew signal input
rlabel metal2 s 537152 -800 537264 480 8 la_data_in[116]
port 180 nsew signal input
rlabel metal2 s 540698 -800 540810 480 8 la_data_in[117]
port 181 nsew signal input
rlabel metal2 s 544244 -800 544356 480 8 la_data_in[118]
port 182 nsew signal input
rlabel metal2 s 547790 -800 547902 480 8 la_data_in[119]
port 183 nsew signal input
rlabel metal2 s 164822 -800 164934 480 8 la_data_in[11]
port 184 nsew signal input
rlabel metal2 s 551336 -800 551448 480 8 la_data_in[120]
port 185 nsew signal input
rlabel metal2 s 554882 -800 554994 480 8 la_data_in[121]
port 186 nsew signal input
rlabel metal2 s 558428 -800 558540 480 8 la_data_in[122]
port 187 nsew signal input
rlabel metal2 s 561974 -800 562086 480 8 la_data_in[123]
port 188 nsew signal input
rlabel metal2 s 565520 -800 565632 480 8 la_data_in[124]
port 189 nsew signal input
rlabel metal2 s 569066 -800 569178 480 8 la_data_in[125]
port 190 nsew signal input
rlabel metal2 s 572612 -800 572724 480 8 la_data_in[126]
port 191 nsew signal input
rlabel metal2 s 576158 -800 576270 480 8 la_data_in[127]
port 192 nsew signal input
rlabel metal2 s 168368 -800 168480 480 8 la_data_in[12]
port 193 nsew signal input
rlabel metal2 s 171914 -800 172026 480 8 la_data_in[13]
port 194 nsew signal input
rlabel metal2 s 175460 -800 175572 480 8 la_data_in[14]
port 195 nsew signal input
rlabel metal2 s 179006 -800 179118 480 8 la_data_in[15]
port 196 nsew signal input
rlabel metal2 s 182552 -800 182664 480 8 la_data_in[16]
port 197 nsew signal input
rlabel metal2 s 186098 -800 186210 480 8 la_data_in[17]
port 198 nsew signal input
rlabel metal2 s 189644 -800 189756 480 8 la_data_in[18]
port 199 nsew signal input
rlabel metal2 s 193190 -800 193302 480 8 la_data_in[19]
port 200 nsew signal input
rlabel metal2 s 129362 -800 129474 480 8 la_data_in[1]
port 201 nsew signal input
rlabel metal2 s 196736 -800 196848 480 8 la_data_in[20]
port 202 nsew signal input
rlabel metal2 s 200282 -800 200394 480 8 la_data_in[21]
port 203 nsew signal input
rlabel metal2 s 203828 -800 203940 480 8 la_data_in[22]
port 204 nsew signal input
rlabel metal2 s 207374 -800 207486 480 8 la_data_in[23]
port 205 nsew signal input
rlabel metal2 s 210920 -800 211032 480 8 la_data_in[24]
port 206 nsew signal input
rlabel metal2 s 214466 -800 214578 480 8 la_data_in[25]
port 207 nsew signal input
rlabel metal2 s 218012 -800 218124 480 8 la_data_in[26]
port 208 nsew signal input
rlabel metal2 s 221558 -800 221670 480 8 la_data_in[27]
port 209 nsew signal input
rlabel metal2 s 225104 -800 225216 480 8 la_data_in[28]
port 210 nsew signal input
rlabel metal2 s 228650 -800 228762 480 8 la_data_in[29]
port 211 nsew signal input
rlabel metal2 s 132908 -800 133020 480 8 la_data_in[2]
port 212 nsew signal input
rlabel metal2 s 232196 -800 232308 480 8 la_data_in[30]
port 213 nsew signal input
rlabel metal2 s 235742 -800 235854 480 8 la_data_in[31]
port 214 nsew signal input
rlabel metal2 s 239288 -800 239400 480 8 la_data_in[32]
port 215 nsew signal input
rlabel metal2 s 242834 -800 242946 480 8 la_data_in[33]
port 216 nsew signal input
rlabel metal2 s 246380 -800 246492 480 8 la_data_in[34]
port 217 nsew signal input
rlabel metal2 s 249926 -800 250038 480 8 la_data_in[35]
port 218 nsew signal input
rlabel metal2 s 253472 -800 253584 480 8 la_data_in[36]
port 219 nsew signal input
rlabel metal2 s 257018 -800 257130 480 8 la_data_in[37]
port 220 nsew signal input
rlabel metal2 s 260564 -800 260676 480 8 la_data_in[38]
port 221 nsew signal input
rlabel metal2 s 264110 -800 264222 480 8 la_data_in[39]
port 222 nsew signal input
rlabel metal2 s 136454 -800 136566 480 8 la_data_in[3]
port 223 nsew signal input
rlabel metal2 s 267656 -800 267768 480 8 la_data_in[40]
port 224 nsew signal input
rlabel metal2 s 271202 -800 271314 480 8 la_data_in[41]
port 225 nsew signal input
rlabel metal2 s 274748 -800 274860 480 8 la_data_in[42]
port 226 nsew signal input
rlabel metal2 s 278294 -800 278406 480 8 la_data_in[43]
port 227 nsew signal input
rlabel metal2 s 281840 -800 281952 480 8 la_data_in[44]
port 228 nsew signal input
rlabel metal2 s 285386 -800 285498 480 8 la_data_in[45]
port 229 nsew signal input
rlabel metal2 s 288932 -800 289044 480 8 la_data_in[46]
port 230 nsew signal input
rlabel metal2 s 292478 -800 292590 480 8 la_data_in[47]
port 231 nsew signal input
rlabel metal2 s 296024 -800 296136 480 8 la_data_in[48]
port 232 nsew signal input
rlabel metal2 s 299570 -800 299682 480 8 la_data_in[49]
port 233 nsew signal input
rlabel metal2 s 140000 -800 140112 480 8 la_data_in[4]
port 234 nsew signal input
rlabel metal2 s 303116 -800 303228 480 8 la_data_in[50]
port 235 nsew signal input
rlabel metal2 s 306662 -800 306774 480 8 la_data_in[51]
port 236 nsew signal input
rlabel metal2 s 310208 -800 310320 480 8 la_data_in[52]
port 237 nsew signal input
rlabel metal2 s 313754 -800 313866 480 8 la_data_in[53]
port 238 nsew signal input
rlabel metal2 s 317300 -800 317412 480 8 la_data_in[54]
port 239 nsew signal input
rlabel metal2 s 320846 -800 320958 480 8 la_data_in[55]
port 240 nsew signal input
rlabel metal2 s 324392 -800 324504 480 8 la_data_in[56]
port 241 nsew signal input
rlabel metal2 s 327938 -800 328050 480 8 la_data_in[57]
port 242 nsew signal input
rlabel metal2 s 331484 -800 331596 480 8 la_data_in[58]
port 243 nsew signal input
rlabel metal2 s 335030 -800 335142 480 8 la_data_in[59]
port 244 nsew signal input
rlabel metal2 s 143546 -800 143658 480 8 la_data_in[5]
port 245 nsew signal input
rlabel metal2 s 338576 -800 338688 480 8 la_data_in[60]
port 246 nsew signal input
rlabel metal2 s 342122 -800 342234 480 8 la_data_in[61]
port 247 nsew signal input
rlabel metal2 s 345668 -800 345780 480 8 la_data_in[62]
port 248 nsew signal input
rlabel metal2 s 349214 -800 349326 480 8 la_data_in[63]
port 249 nsew signal input
rlabel metal2 s 352760 -800 352872 480 8 la_data_in[64]
port 250 nsew signal input
rlabel metal2 s 356306 -800 356418 480 8 la_data_in[65]
port 251 nsew signal input
rlabel metal2 s 359852 -800 359964 480 8 la_data_in[66]
port 252 nsew signal input
rlabel metal2 s 363398 -800 363510 480 8 la_data_in[67]
port 253 nsew signal input
rlabel metal2 s 366944 -800 367056 480 8 la_data_in[68]
port 254 nsew signal input
rlabel metal2 s 370490 -800 370602 480 8 la_data_in[69]
port 255 nsew signal input
rlabel metal2 s 147092 -800 147204 480 8 la_data_in[6]
port 256 nsew signal input
rlabel metal2 s 374036 -800 374148 480 8 la_data_in[70]
port 257 nsew signal input
rlabel metal2 s 377582 -800 377694 480 8 la_data_in[71]
port 258 nsew signal input
rlabel metal2 s 381128 -800 381240 480 8 la_data_in[72]
port 259 nsew signal input
rlabel metal2 s 384674 -800 384786 480 8 la_data_in[73]
port 260 nsew signal input
rlabel metal2 s 388220 -800 388332 480 8 la_data_in[74]
port 261 nsew signal input
rlabel metal2 s 391766 -800 391878 480 8 la_data_in[75]
port 262 nsew signal input
rlabel metal2 s 395312 -800 395424 480 8 la_data_in[76]
port 263 nsew signal input
rlabel metal2 s 398858 -800 398970 480 8 la_data_in[77]
port 264 nsew signal input
rlabel metal2 s 402404 -800 402516 480 8 la_data_in[78]
port 265 nsew signal input
rlabel metal2 s 405950 -800 406062 480 8 la_data_in[79]
port 266 nsew signal input
rlabel metal2 s 150638 -800 150750 480 8 la_data_in[7]
port 267 nsew signal input
rlabel metal2 s 409496 -800 409608 480 8 la_data_in[80]
port 268 nsew signal input
rlabel metal2 s 413042 -800 413154 480 8 la_data_in[81]
port 269 nsew signal input
rlabel metal2 s 416588 -800 416700 480 8 la_data_in[82]
port 270 nsew signal input
rlabel metal2 s 420134 -800 420246 480 8 la_data_in[83]
port 271 nsew signal input
rlabel metal2 s 423680 -800 423792 480 8 la_data_in[84]
port 272 nsew signal input
rlabel metal2 s 427226 -800 427338 480 8 la_data_in[85]
port 273 nsew signal input
rlabel metal2 s 430772 -800 430884 480 8 la_data_in[86]
port 274 nsew signal input
rlabel metal2 s 434318 -800 434430 480 8 la_data_in[87]
port 275 nsew signal input
rlabel metal2 s 437864 -800 437976 480 8 la_data_in[88]
port 276 nsew signal input
rlabel metal2 s 441410 -800 441522 480 8 la_data_in[89]
port 277 nsew signal input
rlabel metal2 s 154184 -800 154296 480 8 la_data_in[8]
port 278 nsew signal input
rlabel metal2 s 444956 -800 445068 480 8 la_data_in[90]
port 279 nsew signal input
rlabel metal2 s 448502 -800 448614 480 8 la_data_in[91]
port 280 nsew signal input
rlabel metal2 s 452048 -800 452160 480 8 la_data_in[92]
port 281 nsew signal input
rlabel metal2 s 455594 -800 455706 480 8 la_data_in[93]
port 282 nsew signal input
rlabel metal2 s 459140 -800 459252 480 8 la_data_in[94]
port 283 nsew signal input
rlabel metal2 s 462686 -800 462798 480 8 la_data_in[95]
port 284 nsew signal input
rlabel metal2 s 466232 -800 466344 480 8 la_data_in[96]
port 285 nsew signal input
rlabel metal2 s 469778 -800 469890 480 8 la_data_in[97]
port 286 nsew signal input
rlabel metal2 s 473324 -800 473436 480 8 la_data_in[98]
port 287 nsew signal input
rlabel metal2 s 476870 -800 476982 480 8 la_data_in[99]
port 288 nsew signal input
rlabel metal2 s 157730 -800 157842 480 8 la_data_in[9]
port 289 nsew signal input
rlabel metal2 s 126998 -800 127110 480 8 la_data_out[0]
port 290 nsew signal output
rlabel metal2 s 481598 -800 481710 480 8 la_data_out[100]
port 291 nsew signal output
rlabel metal2 s 485144 -800 485256 480 8 la_data_out[101]
port 292 nsew signal output
rlabel metal2 s 488690 -800 488802 480 8 la_data_out[102]
port 293 nsew signal output
rlabel metal2 s 492236 -800 492348 480 8 la_data_out[103]
port 294 nsew signal output
rlabel metal2 s 495782 -800 495894 480 8 la_data_out[104]
port 295 nsew signal output
rlabel metal2 s 499328 -800 499440 480 8 la_data_out[105]
port 296 nsew signal output
rlabel metal2 s 502874 -800 502986 480 8 la_data_out[106]
port 297 nsew signal output
rlabel metal2 s 506420 -800 506532 480 8 la_data_out[107]
port 298 nsew signal output
rlabel metal2 s 509966 -800 510078 480 8 la_data_out[108]
port 299 nsew signal output
rlabel metal2 s 513512 -800 513624 480 8 la_data_out[109]
port 300 nsew signal output
rlabel metal2 s 162458 -800 162570 480 8 la_data_out[10]
port 301 nsew signal output
rlabel metal2 s 517058 -800 517170 480 8 la_data_out[110]
port 302 nsew signal output
rlabel metal2 s 520604 -800 520716 480 8 la_data_out[111]
port 303 nsew signal output
rlabel metal2 s 524150 -800 524262 480 8 la_data_out[112]
port 304 nsew signal output
rlabel metal2 s 527696 -800 527808 480 8 la_data_out[113]
port 305 nsew signal output
rlabel metal2 s 531242 -800 531354 480 8 la_data_out[114]
port 306 nsew signal output
rlabel metal2 s 534788 -800 534900 480 8 la_data_out[115]
port 307 nsew signal output
rlabel metal2 s 538334 -800 538446 480 8 la_data_out[116]
port 308 nsew signal output
rlabel metal2 s 541880 -800 541992 480 8 la_data_out[117]
port 309 nsew signal output
rlabel metal2 s 545426 -800 545538 480 8 la_data_out[118]
port 310 nsew signal output
rlabel metal2 s 548972 -800 549084 480 8 la_data_out[119]
port 311 nsew signal output
rlabel metal2 s 166004 -800 166116 480 8 la_data_out[11]
port 312 nsew signal output
rlabel metal2 s 552518 -800 552630 480 8 la_data_out[120]
port 313 nsew signal output
rlabel metal2 s 556064 -800 556176 480 8 la_data_out[121]
port 314 nsew signal output
rlabel metal2 s 559610 -800 559722 480 8 la_data_out[122]
port 315 nsew signal output
rlabel metal2 s 563156 -800 563268 480 8 la_data_out[123]
port 316 nsew signal output
rlabel metal2 s 566702 -800 566814 480 8 la_data_out[124]
port 317 nsew signal output
rlabel metal2 s 570248 -800 570360 480 8 la_data_out[125]
port 318 nsew signal output
rlabel metal2 s 573794 -800 573906 480 8 la_data_out[126]
port 319 nsew signal output
rlabel metal2 s 577340 -800 577452 480 8 la_data_out[127]
port 320 nsew signal output
rlabel metal2 s 169550 -800 169662 480 8 la_data_out[12]
port 321 nsew signal output
rlabel metal2 s 173096 -800 173208 480 8 la_data_out[13]
port 322 nsew signal output
rlabel metal2 s 176642 -800 176754 480 8 la_data_out[14]
port 323 nsew signal output
rlabel metal2 s 180188 -800 180300 480 8 la_data_out[15]
port 324 nsew signal output
rlabel metal2 s 183734 -800 183846 480 8 la_data_out[16]
port 325 nsew signal output
rlabel metal2 s 187280 -800 187392 480 8 la_data_out[17]
port 326 nsew signal output
rlabel metal2 s 190826 -800 190938 480 8 la_data_out[18]
port 327 nsew signal output
rlabel metal2 s 194372 -800 194484 480 8 la_data_out[19]
port 328 nsew signal output
rlabel metal2 s 130544 -800 130656 480 8 la_data_out[1]
port 329 nsew signal output
rlabel metal2 s 197918 -800 198030 480 8 la_data_out[20]
port 330 nsew signal output
rlabel metal2 s 201464 -800 201576 480 8 la_data_out[21]
port 331 nsew signal output
rlabel metal2 s 205010 -800 205122 480 8 la_data_out[22]
port 332 nsew signal output
rlabel metal2 s 208556 -800 208668 480 8 la_data_out[23]
port 333 nsew signal output
rlabel metal2 s 212102 -800 212214 480 8 la_data_out[24]
port 334 nsew signal output
rlabel metal2 s 215648 -800 215760 480 8 la_data_out[25]
port 335 nsew signal output
rlabel metal2 s 219194 -800 219306 480 8 la_data_out[26]
port 336 nsew signal output
rlabel metal2 s 222740 -800 222852 480 8 la_data_out[27]
port 337 nsew signal output
rlabel metal2 s 226286 -800 226398 480 8 la_data_out[28]
port 338 nsew signal output
rlabel metal2 s 229832 -800 229944 480 8 la_data_out[29]
port 339 nsew signal output
rlabel metal2 s 134090 -800 134202 480 8 la_data_out[2]
port 340 nsew signal output
rlabel metal2 s 233378 -800 233490 480 8 la_data_out[30]
port 341 nsew signal output
rlabel metal2 s 236924 -800 237036 480 8 la_data_out[31]
port 342 nsew signal output
rlabel metal2 s 240470 -800 240582 480 8 la_data_out[32]
port 343 nsew signal output
rlabel metal2 s 244016 -800 244128 480 8 la_data_out[33]
port 344 nsew signal output
rlabel metal2 s 247562 -800 247674 480 8 la_data_out[34]
port 345 nsew signal output
rlabel metal2 s 251108 -800 251220 480 8 la_data_out[35]
port 346 nsew signal output
rlabel metal2 s 254654 -800 254766 480 8 la_data_out[36]
port 347 nsew signal output
rlabel metal2 s 258200 -800 258312 480 8 la_data_out[37]
port 348 nsew signal output
rlabel metal2 s 261746 -800 261858 480 8 la_data_out[38]
port 349 nsew signal output
rlabel metal2 s 265292 -800 265404 480 8 la_data_out[39]
port 350 nsew signal output
rlabel metal2 s 137636 -800 137748 480 8 la_data_out[3]
port 351 nsew signal output
rlabel metal2 s 268838 -800 268950 480 8 la_data_out[40]
port 352 nsew signal output
rlabel metal2 s 272384 -800 272496 480 8 la_data_out[41]
port 353 nsew signal output
rlabel metal2 s 275930 -800 276042 480 8 la_data_out[42]
port 354 nsew signal output
rlabel metal2 s 279476 -800 279588 480 8 la_data_out[43]
port 355 nsew signal output
rlabel metal2 s 283022 -800 283134 480 8 la_data_out[44]
port 356 nsew signal output
rlabel metal2 s 286568 -800 286680 480 8 la_data_out[45]
port 357 nsew signal output
rlabel metal2 s 290114 -800 290226 480 8 la_data_out[46]
port 358 nsew signal output
rlabel metal2 s 293660 -800 293772 480 8 la_data_out[47]
port 359 nsew signal output
rlabel metal2 s 297206 -800 297318 480 8 la_data_out[48]
port 360 nsew signal output
rlabel metal2 s 300752 -800 300864 480 8 la_data_out[49]
port 361 nsew signal output
rlabel metal2 s 141182 -800 141294 480 8 la_data_out[4]
port 362 nsew signal output
rlabel metal2 s 304298 -800 304410 480 8 la_data_out[50]
port 363 nsew signal output
rlabel metal2 s 307844 -800 307956 480 8 la_data_out[51]
port 364 nsew signal output
rlabel metal2 s 311390 -800 311502 480 8 la_data_out[52]
port 365 nsew signal output
rlabel metal2 s 314936 -800 315048 480 8 la_data_out[53]
port 366 nsew signal output
rlabel metal2 s 318482 -800 318594 480 8 la_data_out[54]
port 367 nsew signal output
rlabel metal2 s 322028 -800 322140 480 8 la_data_out[55]
port 368 nsew signal output
rlabel metal2 s 325574 -800 325686 480 8 la_data_out[56]
port 369 nsew signal output
rlabel metal2 s 329120 -800 329232 480 8 la_data_out[57]
port 370 nsew signal output
rlabel metal2 s 332666 -800 332778 480 8 la_data_out[58]
port 371 nsew signal output
rlabel metal2 s 336212 -800 336324 480 8 la_data_out[59]
port 372 nsew signal output
rlabel metal2 s 144728 -800 144840 480 8 la_data_out[5]
port 373 nsew signal output
rlabel metal2 s 339758 -800 339870 480 8 la_data_out[60]
port 374 nsew signal output
rlabel metal2 s 343304 -800 343416 480 8 la_data_out[61]
port 375 nsew signal output
rlabel metal2 s 346850 -800 346962 480 8 la_data_out[62]
port 376 nsew signal output
rlabel metal2 s 350396 -800 350508 480 8 la_data_out[63]
port 377 nsew signal output
rlabel metal2 s 353942 -800 354054 480 8 la_data_out[64]
port 378 nsew signal output
rlabel metal2 s 357488 -800 357600 480 8 la_data_out[65]
port 379 nsew signal output
rlabel metal2 s 361034 -800 361146 480 8 la_data_out[66]
port 380 nsew signal output
rlabel metal2 s 364580 -800 364692 480 8 la_data_out[67]
port 381 nsew signal output
rlabel metal2 s 368126 -800 368238 480 8 la_data_out[68]
port 382 nsew signal output
rlabel metal2 s 371672 -800 371784 480 8 la_data_out[69]
port 383 nsew signal output
rlabel metal2 s 148274 -800 148386 480 8 la_data_out[6]
port 384 nsew signal output
rlabel metal2 s 375218 -800 375330 480 8 la_data_out[70]
port 385 nsew signal output
rlabel metal2 s 378764 -800 378876 480 8 la_data_out[71]
port 386 nsew signal output
rlabel metal2 s 382310 -800 382422 480 8 la_data_out[72]
port 387 nsew signal output
rlabel metal2 s 385856 -800 385968 480 8 la_data_out[73]
port 388 nsew signal output
rlabel metal2 s 389402 -800 389514 480 8 la_data_out[74]
port 389 nsew signal output
rlabel metal2 s 392948 -800 393060 480 8 la_data_out[75]
port 390 nsew signal output
rlabel metal2 s 396494 -800 396606 480 8 la_data_out[76]
port 391 nsew signal output
rlabel metal2 s 400040 -800 400152 480 8 la_data_out[77]
port 392 nsew signal output
rlabel metal2 s 403586 -800 403698 480 8 la_data_out[78]
port 393 nsew signal output
rlabel metal2 s 407132 -800 407244 480 8 la_data_out[79]
port 394 nsew signal output
rlabel metal2 s 151820 -800 151932 480 8 la_data_out[7]
port 395 nsew signal output
rlabel metal2 s 410678 -800 410790 480 8 la_data_out[80]
port 396 nsew signal output
rlabel metal2 s 414224 -800 414336 480 8 la_data_out[81]
port 397 nsew signal output
rlabel metal2 s 417770 -800 417882 480 8 la_data_out[82]
port 398 nsew signal output
rlabel metal2 s 421316 -800 421428 480 8 la_data_out[83]
port 399 nsew signal output
rlabel metal2 s 424862 -800 424974 480 8 la_data_out[84]
port 400 nsew signal output
rlabel metal2 s 428408 -800 428520 480 8 la_data_out[85]
port 401 nsew signal output
rlabel metal2 s 431954 -800 432066 480 8 la_data_out[86]
port 402 nsew signal output
rlabel metal2 s 435500 -800 435612 480 8 la_data_out[87]
port 403 nsew signal output
rlabel metal2 s 439046 -800 439158 480 8 la_data_out[88]
port 404 nsew signal output
rlabel metal2 s 442592 -800 442704 480 8 la_data_out[89]
port 405 nsew signal output
rlabel metal2 s 155366 -800 155478 480 8 la_data_out[8]
port 406 nsew signal output
rlabel metal2 s 446138 -800 446250 480 8 la_data_out[90]
port 407 nsew signal output
rlabel metal2 s 449684 -800 449796 480 8 la_data_out[91]
port 408 nsew signal output
rlabel metal2 s 453230 -800 453342 480 8 la_data_out[92]
port 409 nsew signal output
rlabel metal2 s 456776 -800 456888 480 8 la_data_out[93]
port 410 nsew signal output
rlabel metal2 s 460322 -800 460434 480 8 la_data_out[94]
port 411 nsew signal output
rlabel metal2 s 463868 -800 463980 480 8 la_data_out[95]
port 412 nsew signal output
rlabel metal2 s 467414 -800 467526 480 8 la_data_out[96]
port 413 nsew signal output
rlabel metal2 s 470960 -800 471072 480 8 la_data_out[97]
port 414 nsew signal output
rlabel metal2 s 474506 -800 474618 480 8 la_data_out[98]
port 415 nsew signal output
rlabel metal2 s 478052 -800 478164 480 8 la_data_out[99]
port 416 nsew signal output
rlabel metal2 s 158912 -800 159024 480 8 la_data_out[9]
port 417 nsew signal output
rlabel metal2 s 128180 -800 128292 480 8 la_oenb[0]
port 418 nsew signal input
rlabel metal2 s 482780 -800 482892 480 8 la_oenb[100]
port 419 nsew signal input
rlabel metal2 s 486326 -800 486438 480 8 la_oenb[101]
port 420 nsew signal input
rlabel metal2 s 489872 -800 489984 480 8 la_oenb[102]
port 421 nsew signal input
rlabel metal2 s 493418 -800 493530 480 8 la_oenb[103]
port 422 nsew signal input
rlabel metal2 s 496964 -800 497076 480 8 la_oenb[104]
port 423 nsew signal input
rlabel metal2 s 500510 -800 500622 480 8 la_oenb[105]
port 424 nsew signal input
rlabel metal2 s 504056 -800 504168 480 8 la_oenb[106]
port 425 nsew signal input
rlabel metal2 s 507602 -800 507714 480 8 la_oenb[107]
port 426 nsew signal input
rlabel metal2 s 511148 -800 511260 480 8 la_oenb[108]
port 427 nsew signal input
rlabel metal2 s 514694 -800 514806 480 8 la_oenb[109]
port 428 nsew signal input
rlabel metal2 s 163640 -800 163752 480 8 la_oenb[10]
port 429 nsew signal input
rlabel metal2 s 518240 -800 518352 480 8 la_oenb[110]
port 430 nsew signal input
rlabel metal2 s 521786 -800 521898 480 8 la_oenb[111]
port 431 nsew signal input
rlabel metal2 s 525332 -800 525444 480 8 la_oenb[112]
port 432 nsew signal input
rlabel metal2 s 528878 -800 528990 480 8 la_oenb[113]
port 433 nsew signal input
rlabel metal2 s 532424 -800 532536 480 8 la_oenb[114]
port 434 nsew signal input
rlabel metal2 s 535970 -800 536082 480 8 la_oenb[115]
port 435 nsew signal input
rlabel metal2 s 539516 -800 539628 480 8 la_oenb[116]
port 436 nsew signal input
rlabel metal2 s 543062 -800 543174 480 8 la_oenb[117]
port 437 nsew signal input
rlabel metal2 s 546608 -800 546720 480 8 la_oenb[118]
port 438 nsew signal input
rlabel metal2 s 550154 -800 550266 480 8 la_oenb[119]
port 439 nsew signal input
rlabel metal2 s 167186 -800 167298 480 8 la_oenb[11]
port 440 nsew signal input
rlabel metal2 s 553700 -800 553812 480 8 la_oenb[120]
port 441 nsew signal input
rlabel metal2 s 557246 -800 557358 480 8 la_oenb[121]
port 442 nsew signal input
rlabel metal2 s 560792 -800 560904 480 8 la_oenb[122]
port 443 nsew signal input
rlabel metal2 s 564338 -800 564450 480 8 la_oenb[123]
port 444 nsew signal input
rlabel metal2 s 567884 -800 567996 480 8 la_oenb[124]
port 445 nsew signal input
rlabel metal2 s 571430 -800 571542 480 8 la_oenb[125]
port 446 nsew signal input
rlabel metal2 s 574976 -800 575088 480 8 la_oenb[126]
port 447 nsew signal input
rlabel metal2 s 578522 -800 578634 480 8 la_oenb[127]
port 448 nsew signal input
rlabel metal2 s 170732 -800 170844 480 8 la_oenb[12]
port 449 nsew signal input
rlabel metal2 s 174278 -800 174390 480 8 la_oenb[13]
port 450 nsew signal input
rlabel metal2 s 177824 -800 177936 480 8 la_oenb[14]
port 451 nsew signal input
rlabel metal2 s 181370 -800 181482 480 8 la_oenb[15]
port 452 nsew signal input
rlabel metal2 s 184916 -800 185028 480 8 la_oenb[16]
port 453 nsew signal input
rlabel metal2 s 188462 -800 188574 480 8 la_oenb[17]
port 454 nsew signal input
rlabel metal2 s 192008 -800 192120 480 8 la_oenb[18]
port 455 nsew signal input
rlabel metal2 s 195554 -800 195666 480 8 la_oenb[19]
port 456 nsew signal input
rlabel metal2 s 131726 -800 131838 480 8 la_oenb[1]
port 457 nsew signal input
rlabel metal2 s 199100 -800 199212 480 8 la_oenb[20]
port 458 nsew signal input
rlabel metal2 s 202646 -800 202758 480 8 la_oenb[21]
port 459 nsew signal input
rlabel metal2 s 206192 -800 206304 480 8 la_oenb[22]
port 460 nsew signal input
rlabel metal2 s 209738 -800 209850 480 8 la_oenb[23]
port 461 nsew signal input
rlabel metal2 s 213284 -800 213396 480 8 la_oenb[24]
port 462 nsew signal input
rlabel metal2 s 216830 -800 216942 480 8 la_oenb[25]
port 463 nsew signal input
rlabel metal2 s 220376 -800 220488 480 8 la_oenb[26]
port 464 nsew signal input
rlabel metal2 s 223922 -800 224034 480 8 la_oenb[27]
port 465 nsew signal input
rlabel metal2 s 227468 -800 227580 480 8 la_oenb[28]
port 466 nsew signal input
rlabel metal2 s 231014 -800 231126 480 8 la_oenb[29]
port 467 nsew signal input
rlabel metal2 s 135272 -800 135384 480 8 la_oenb[2]
port 468 nsew signal input
rlabel metal2 s 234560 -800 234672 480 8 la_oenb[30]
port 469 nsew signal input
rlabel metal2 s 238106 -800 238218 480 8 la_oenb[31]
port 470 nsew signal input
rlabel metal2 s 241652 -800 241764 480 8 la_oenb[32]
port 471 nsew signal input
rlabel metal2 s 245198 -800 245310 480 8 la_oenb[33]
port 472 nsew signal input
rlabel metal2 s 248744 -800 248856 480 8 la_oenb[34]
port 473 nsew signal input
rlabel metal2 s 252290 -800 252402 480 8 la_oenb[35]
port 474 nsew signal input
rlabel metal2 s 255836 -800 255948 480 8 la_oenb[36]
port 475 nsew signal input
rlabel metal2 s 259382 -800 259494 480 8 la_oenb[37]
port 476 nsew signal input
rlabel metal2 s 262928 -800 263040 480 8 la_oenb[38]
port 477 nsew signal input
rlabel metal2 s 266474 -800 266586 480 8 la_oenb[39]
port 478 nsew signal input
rlabel metal2 s 138818 -800 138930 480 8 la_oenb[3]
port 479 nsew signal input
rlabel metal2 s 270020 -800 270132 480 8 la_oenb[40]
port 480 nsew signal input
rlabel metal2 s 273566 -800 273678 480 8 la_oenb[41]
port 481 nsew signal input
rlabel metal2 s 277112 -800 277224 480 8 la_oenb[42]
port 482 nsew signal input
rlabel metal2 s 280658 -800 280770 480 8 la_oenb[43]
port 483 nsew signal input
rlabel metal2 s 284204 -800 284316 480 8 la_oenb[44]
port 484 nsew signal input
rlabel metal2 s 287750 -800 287862 480 8 la_oenb[45]
port 485 nsew signal input
rlabel metal2 s 291296 -800 291408 480 8 la_oenb[46]
port 486 nsew signal input
rlabel metal2 s 294842 -800 294954 480 8 la_oenb[47]
port 487 nsew signal input
rlabel metal2 s 298388 -800 298500 480 8 la_oenb[48]
port 488 nsew signal input
rlabel metal2 s 301934 -800 302046 480 8 la_oenb[49]
port 489 nsew signal input
rlabel metal2 s 142364 -800 142476 480 8 la_oenb[4]
port 490 nsew signal input
rlabel metal2 s 305480 -800 305592 480 8 la_oenb[50]
port 491 nsew signal input
rlabel metal2 s 309026 -800 309138 480 8 la_oenb[51]
port 492 nsew signal input
rlabel metal2 s 312572 -800 312684 480 8 la_oenb[52]
port 493 nsew signal input
rlabel metal2 s 316118 -800 316230 480 8 la_oenb[53]
port 494 nsew signal input
rlabel metal2 s 319664 -800 319776 480 8 la_oenb[54]
port 495 nsew signal input
rlabel metal2 s 323210 -800 323322 480 8 la_oenb[55]
port 496 nsew signal input
rlabel metal2 s 326756 -800 326868 480 8 la_oenb[56]
port 497 nsew signal input
rlabel metal2 s 330302 -800 330414 480 8 la_oenb[57]
port 498 nsew signal input
rlabel metal2 s 333848 -800 333960 480 8 la_oenb[58]
port 499 nsew signal input
rlabel metal2 s 337394 -800 337506 480 8 la_oenb[59]
port 500 nsew signal input
rlabel metal2 s 145910 -800 146022 480 8 la_oenb[5]
port 501 nsew signal input
rlabel metal2 s 340940 -800 341052 480 8 la_oenb[60]
port 502 nsew signal input
rlabel metal2 s 344486 -800 344598 480 8 la_oenb[61]
port 503 nsew signal input
rlabel metal2 s 348032 -800 348144 480 8 la_oenb[62]
port 504 nsew signal input
rlabel metal2 s 351578 -800 351690 480 8 la_oenb[63]
port 505 nsew signal input
rlabel metal2 s 355124 -800 355236 480 8 la_oenb[64]
port 506 nsew signal input
rlabel metal2 s 358670 -800 358782 480 8 la_oenb[65]
port 507 nsew signal input
rlabel metal2 s 362216 -800 362328 480 8 la_oenb[66]
port 508 nsew signal input
rlabel metal2 s 365762 -800 365874 480 8 la_oenb[67]
port 509 nsew signal input
rlabel metal2 s 369308 -800 369420 480 8 la_oenb[68]
port 510 nsew signal input
rlabel metal2 s 372854 -800 372966 480 8 la_oenb[69]
port 511 nsew signal input
rlabel metal2 s 149456 -800 149568 480 8 la_oenb[6]
port 512 nsew signal input
rlabel metal2 s 376400 -800 376512 480 8 la_oenb[70]
port 513 nsew signal input
rlabel metal2 s 379946 -800 380058 480 8 la_oenb[71]
port 514 nsew signal input
rlabel metal2 s 383492 -800 383604 480 8 la_oenb[72]
port 515 nsew signal input
rlabel metal2 s 387038 -800 387150 480 8 la_oenb[73]
port 516 nsew signal input
rlabel metal2 s 390584 -800 390696 480 8 la_oenb[74]
port 517 nsew signal input
rlabel metal2 s 394130 -800 394242 480 8 la_oenb[75]
port 518 nsew signal input
rlabel metal2 s 397676 -800 397788 480 8 la_oenb[76]
port 519 nsew signal input
rlabel metal2 s 401222 -800 401334 480 8 la_oenb[77]
port 520 nsew signal input
rlabel metal2 s 404768 -800 404880 480 8 la_oenb[78]
port 521 nsew signal input
rlabel metal2 s 408314 -800 408426 480 8 la_oenb[79]
port 522 nsew signal input
rlabel metal2 s 153002 -800 153114 480 8 la_oenb[7]
port 523 nsew signal input
rlabel metal2 s 411860 -800 411972 480 8 la_oenb[80]
port 524 nsew signal input
rlabel metal2 s 415406 -800 415518 480 8 la_oenb[81]
port 525 nsew signal input
rlabel metal2 s 418952 -800 419064 480 8 la_oenb[82]
port 526 nsew signal input
rlabel metal2 s 422498 -800 422610 480 8 la_oenb[83]
port 527 nsew signal input
rlabel metal2 s 426044 -800 426156 480 8 la_oenb[84]
port 528 nsew signal input
rlabel metal2 s 429590 -800 429702 480 8 la_oenb[85]
port 529 nsew signal input
rlabel metal2 s 433136 -800 433248 480 8 la_oenb[86]
port 530 nsew signal input
rlabel metal2 s 436682 -800 436794 480 8 la_oenb[87]
port 531 nsew signal input
rlabel metal2 s 440228 -800 440340 480 8 la_oenb[88]
port 532 nsew signal input
rlabel metal2 s 443774 -800 443886 480 8 la_oenb[89]
port 533 nsew signal input
rlabel metal2 s 156548 -800 156660 480 8 la_oenb[8]
port 534 nsew signal input
rlabel metal2 s 447320 -800 447432 480 8 la_oenb[90]
port 535 nsew signal input
rlabel metal2 s 450866 -800 450978 480 8 la_oenb[91]
port 536 nsew signal input
rlabel metal2 s 454412 -800 454524 480 8 la_oenb[92]
port 537 nsew signal input
rlabel metal2 s 457958 -800 458070 480 8 la_oenb[93]
port 538 nsew signal input
rlabel metal2 s 461504 -800 461616 480 8 la_oenb[94]
port 539 nsew signal input
rlabel metal2 s 465050 -800 465162 480 8 la_oenb[95]
port 540 nsew signal input
rlabel metal2 s 468596 -800 468708 480 8 la_oenb[96]
port 541 nsew signal input
rlabel metal2 s 472142 -800 472254 480 8 la_oenb[97]
port 542 nsew signal input
rlabel metal2 s 475688 -800 475800 480 8 la_oenb[98]
port 543 nsew signal input
rlabel metal2 s 479234 -800 479346 480 8 la_oenb[99]
port 544 nsew signal input
rlabel metal2 s 160094 -800 160206 480 8 la_oenb[9]
port 545 nsew signal input
rlabel metal2 s 579704 -800 579816 480 8 user_clock2
port 546 nsew signal input
rlabel metal2 s 580886 -800 580998 480 8 user_irq[0]
port 547 nsew signal output
rlabel metal2 s 582068 -800 582180 480 8 user_irq[1]
port 548 nsew signal output
rlabel metal2 s 583250 -800 583362 480 8 user_irq[2]
port 549 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 550 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 550 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 9234 -7654 9854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 45234 -7654 45854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 81234 -7654 81854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 117234 -7654 117854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 153234 -7654 153854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 189234 -7654 189854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 225234 -7654 225854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 261234 102564 261854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 297234 -7654 297854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 333234 -7654 333854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 369234 102564 369854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 405234 -7654 405854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 441234 -7654 441854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 477234 102564 477854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 513234 -7654 513854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s 549234 -7654 549854 711590 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 10306 592650 10926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 46306 592650 46926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 82306 592650 82926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 118306 592650 118926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 154306 592650 154926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 190306 592650 190926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 226306 592650 226926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 262306 592650 262926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 298306 592650 298926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 334306 592650 334926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 370306 592650 370926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 406306 592650 406926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 442306 592650 442926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 478306 592650 478926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 514306 592650 514926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 550306 592650 550926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 586306 592650 586926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 622306 592650 622926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 658306 592650 658926 6 vccd2
port 551 nsew power bidirectional
rlabel metal5 s -8726 694306 592650 694926 6 vccd2
port 551 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 16674 -7654 17294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 52674 -7654 53294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 88674 -7654 89294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 124674 -7654 125294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 160674 -7654 161294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 196674 -7654 197294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 232674 -7654 233294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 268674 -7654 269294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 304674 -7654 305294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 340674 -7654 341294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 376674 -7654 377294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 412674 -7654 413294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 448674 -7654 449294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 484674 -7654 485294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 520674 -7654 521294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s 556674 -7654 557294 711590 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 17746 592650 18366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 53746 592650 54366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 89746 592650 90366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 125746 592650 126366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 161746 592650 162366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 197746 592650 198366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 233746 592650 234366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 269746 592650 270366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 305746 592650 306366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 341746 592650 342366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 377746 592650 378366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 413746 592650 414366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 449746 592650 450366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 485746 592650 486366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 521746 592650 522366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 557746 592650 558366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 593746 592650 594366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 629746 592650 630366 6 vdda1
port 552 nsew power bidirectional
rlabel metal5 s -8726 665746 592650 666366 6 vdda1
port 552 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 24114 -7654 24734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 60114 -7654 60734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 96114 -7654 96734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 132114 -7654 132734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 168114 -7654 168734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 204114 -7654 204734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 240114 -7654 240734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 276114 -7654 276734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 312114 -7654 312734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 348114 -7654 348734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 384114 102564 384734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 420114 -7654 420734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 456114 -7654 456734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 492114 102564 492734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 528114 -7654 528734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s 564114 -7654 564734 711590 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 25186 592650 25806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 61186 592650 61806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 97186 592650 97806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 133186 592650 133806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 169186 592650 169806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 205186 592650 205806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 241186 592650 241806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 277186 592650 277806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 313186 592650 313806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 349186 592650 349806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 385186 592650 385806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 421186 592650 421806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 457186 592650 457806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 493186 592650 493806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 529186 592650 529806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 565186 592650 565806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 601186 592650 601806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 637186 592650 637806 6 vdda2
port 553 nsew power bidirectional
rlabel metal5 s -8726 673186 592650 673806 6 vdda2
port 553 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 20394 -7654 21014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 56394 -7654 57014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 92394 102564 93014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 128394 -7654 129014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 164394 -7654 165014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 200394 102564 201014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 236394 -7654 237014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 272394 -7654 273014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 308394 102564 309014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 344394 -7654 345014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 380394 -7654 381014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 416394 -7654 417014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 452394 -7654 453014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 488394 -7654 489014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 524394 -7654 525014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s 560394 -7654 561014 711590 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 21466 592650 22086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 57466 592650 58086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 93466 592650 94086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 129466 592650 130086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 165466 592650 166086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 201466 592650 202086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 237466 592650 238086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 273466 592650 274086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 309466 592650 310086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 345466 592650 346086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 381466 592650 382086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 417466 592650 418086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 453466 592650 454086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 489466 592650 490086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 525466 592650 526086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 561466 592650 562086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 597466 592650 598086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 633466 592650 634086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal5 s -8726 669466 592650 670086 6 vssa1
port 554 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 27834 -7654 28454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 63834 -7654 64454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 99834 -7654 100454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 135834 -7654 136454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 171834 -7654 172454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 207834 -7654 208454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 243834 -7654 244454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 279834 -7654 280454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 315834 -7654 316454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 351834 -7654 352454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 387834 -7654 388454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 423834 -7654 424454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 459834 -7654 460454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 495834 -7654 496454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 531834 -7654 532454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s 567834 -7654 568454 711590 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 28906 592650 29526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 64906 592650 65526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 100906 592650 101526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 136906 592650 137526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 172906 592650 173526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 208906 592650 209526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 244906 592650 245526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 280906 592650 281526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 316906 592650 317526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 352906 592650 353526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 388906 592650 389526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 424906 592650 425526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 460906 592650 461526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 496906 592650 497526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 532906 592650 533526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 568906 592650 569526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 604906 592650 605526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 640906 592650 641526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal5 s -8726 676906 592650 677526 6 vssa2
port 555 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 5514 -7654 6134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 41514 -7654 42134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 77514 102564 78134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 113514 -7654 114134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 149514 -7654 150134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 185514 102564 186134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 221514 -7654 222134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 257514 -7654 258134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 293514 -7654 294134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 329514 -7654 330134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 365514 -7654 366134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 401514 -7654 402134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 437514 -7654 438134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 473514 -7654 474134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 509514 -7654 510134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 545514 -7654 546134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s 581514 -7654 582134 711590 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 6586 592650 7206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 42586 592650 43206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 78586 592650 79206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 114586 592650 115206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 150586 592650 151206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 186586 592650 187206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 222586 592650 223206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 258586 592650 259206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 294586 592650 295206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 330586 592650 331206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 366586 592650 367206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 402586 592650 403206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 438586 592650 439206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 474586 592650 475206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 510586 592650 511206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 546586 592650 547206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 582586 592650 583206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 618586 592650 619206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 654586 592650 655206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal5 s -8726 690586 592650 691206 6 vssd1
port 556 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 12954 -7654 13574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 48954 -7654 49574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 84954 -7654 85574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 120954 -7654 121574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 156954 -7654 157574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 192954 -7654 193574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 228954 -7654 229574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 264954 -7654 265574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 300954 -7654 301574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 336954 -7654 337574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 372954 -7654 373574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 408954 -7654 409574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 444954 -7654 445574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 480954 -7654 481574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 516954 -7654 517574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal4 s 552954 -7654 553574 711590 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 14026 592650 14646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 50026 592650 50646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 86026 592650 86646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 122026 592650 122646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 158026 592650 158646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 194026 592650 194646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 230026 592650 230646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 266026 592650 266646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 302026 592650 302646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 338026 592650 338646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 374026 592650 374646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 410026 592650 410646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 446026 592650 446646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 482026 592650 482646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 518026 592650 518646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 554026 592650 554646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 590026 592650 590646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 626026 592650 626646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 662026 592650 662646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal5 s -8726 698026 592650 698646 6 vssd2
port 557 nsew ground bidirectional
rlabel metal2 s 524 -800 636 480 8 wb_clk_i
port 558 nsew signal input
rlabel metal2 s 1706 -800 1818 480 8 wb_rst_i
port 559 nsew signal input
rlabel metal2 s 2888 -800 3000 480 8 wbs_ack_o
port 560 nsew signal output
rlabel metal2 s 7616 -800 7728 480 8 wbs_adr_i[0]
port 561 nsew signal input
rlabel metal2 s 47804 -800 47916 480 8 wbs_adr_i[10]
port 562 nsew signal input
rlabel metal2 s 51350 -800 51462 480 8 wbs_adr_i[11]
port 563 nsew signal input
rlabel metal2 s 54896 -800 55008 480 8 wbs_adr_i[12]
port 564 nsew signal input
rlabel metal2 s 58442 -800 58554 480 8 wbs_adr_i[13]
port 565 nsew signal input
rlabel metal2 s 61988 -800 62100 480 8 wbs_adr_i[14]
port 566 nsew signal input
rlabel metal2 s 65534 -800 65646 480 8 wbs_adr_i[15]
port 567 nsew signal input
rlabel metal2 s 69080 -800 69192 480 8 wbs_adr_i[16]
port 568 nsew signal input
rlabel metal2 s 72626 -800 72738 480 8 wbs_adr_i[17]
port 569 nsew signal input
rlabel metal2 s 76172 -800 76284 480 8 wbs_adr_i[18]
port 570 nsew signal input
rlabel metal2 s 79718 -800 79830 480 8 wbs_adr_i[19]
port 571 nsew signal input
rlabel metal2 s 12344 -800 12456 480 8 wbs_adr_i[1]
port 572 nsew signal input
rlabel metal2 s 83264 -800 83376 480 8 wbs_adr_i[20]
port 573 nsew signal input
rlabel metal2 s 86810 -800 86922 480 8 wbs_adr_i[21]
port 574 nsew signal input
rlabel metal2 s 90356 -800 90468 480 8 wbs_adr_i[22]
port 575 nsew signal input
rlabel metal2 s 93902 -800 94014 480 8 wbs_adr_i[23]
port 576 nsew signal input
rlabel metal2 s 97448 -800 97560 480 8 wbs_adr_i[24]
port 577 nsew signal input
rlabel metal2 s 100994 -800 101106 480 8 wbs_adr_i[25]
port 578 nsew signal input
rlabel metal2 s 104540 -800 104652 480 8 wbs_adr_i[26]
port 579 nsew signal input
rlabel metal2 s 108086 -800 108198 480 8 wbs_adr_i[27]
port 580 nsew signal input
rlabel metal2 s 111632 -800 111744 480 8 wbs_adr_i[28]
port 581 nsew signal input
rlabel metal2 s 115178 -800 115290 480 8 wbs_adr_i[29]
port 582 nsew signal input
rlabel metal2 s 17072 -800 17184 480 8 wbs_adr_i[2]
port 583 nsew signal input
rlabel metal2 s 118724 -800 118836 480 8 wbs_adr_i[30]
port 584 nsew signal input
rlabel metal2 s 122270 -800 122382 480 8 wbs_adr_i[31]
port 585 nsew signal input
rlabel metal2 s 21800 -800 21912 480 8 wbs_adr_i[3]
port 586 nsew signal input
rlabel metal2 s 26528 -800 26640 480 8 wbs_adr_i[4]
port 587 nsew signal input
rlabel metal2 s 30074 -800 30186 480 8 wbs_adr_i[5]
port 588 nsew signal input
rlabel metal2 s 33620 -800 33732 480 8 wbs_adr_i[6]
port 589 nsew signal input
rlabel metal2 s 37166 -800 37278 480 8 wbs_adr_i[7]
port 590 nsew signal input
rlabel metal2 s 40712 -800 40824 480 8 wbs_adr_i[8]
port 591 nsew signal input
rlabel metal2 s 44258 -800 44370 480 8 wbs_adr_i[9]
port 592 nsew signal input
rlabel metal2 s 4070 -800 4182 480 8 wbs_cyc_i
port 593 nsew signal input
rlabel metal2 s 8798 -800 8910 480 8 wbs_dat_i[0]
port 594 nsew signal input
rlabel metal2 s 48986 -800 49098 480 8 wbs_dat_i[10]
port 595 nsew signal input
rlabel metal2 s 52532 -800 52644 480 8 wbs_dat_i[11]
port 596 nsew signal input
rlabel metal2 s 56078 -800 56190 480 8 wbs_dat_i[12]
port 597 nsew signal input
rlabel metal2 s 59624 -800 59736 480 8 wbs_dat_i[13]
port 598 nsew signal input
rlabel metal2 s 63170 -800 63282 480 8 wbs_dat_i[14]
port 599 nsew signal input
rlabel metal2 s 66716 -800 66828 480 8 wbs_dat_i[15]
port 600 nsew signal input
rlabel metal2 s 70262 -800 70374 480 8 wbs_dat_i[16]
port 601 nsew signal input
rlabel metal2 s 73808 -800 73920 480 8 wbs_dat_i[17]
port 602 nsew signal input
rlabel metal2 s 77354 -800 77466 480 8 wbs_dat_i[18]
port 603 nsew signal input
rlabel metal2 s 80900 -800 81012 480 8 wbs_dat_i[19]
port 604 nsew signal input
rlabel metal2 s 13526 -800 13638 480 8 wbs_dat_i[1]
port 605 nsew signal input
rlabel metal2 s 84446 -800 84558 480 8 wbs_dat_i[20]
port 606 nsew signal input
rlabel metal2 s 87992 -800 88104 480 8 wbs_dat_i[21]
port 607 nsew signal input
rlabel metal2 s 91538 -800 91650 480 8 wbs_dat_i[22]
port 608 nsew signal input
rlabel metal2 s 95084 -800 95196 480 8 wbs_dat_i[23]
port 609 nsew signal input
rlabel metal2 s 98630 -800 98742 480 8 wbs_dat_i[24]
port 610 nsew signal input
rlabel metal2 s 102176 -800 102288 480 8 wbs_dat_i[25]
port 611 nsew signal input
rlabel metal2 s 105722 -800 105834 480 8 wbs_dat_i[26]
port 612 nsew signal input
rlabel metal2 s 109268 -800 109380 480 8 wbs_dat_i[27]
port 613 nsew signal input
rlabel metal2 s 112814 -800 112926 480 8 wbs_dat_i[28]
port 614 nsew signal input
rlabel metal2 s 116360 -800 116472 480 8 wbs_dat_i[29]
port 615 nsew signal input
rlabel metal2 s 18254 -800 18366 480 8 wbs_dat_i[2]
port 616 nsew signal input
rlabel metal2 s 119906 -800 120018 480 8 wbs_dat_i[30]
port 617 nsew signal input
rlabel metal2 s 123452 -800 123564 480 8 wbs_dat_i[31]
port 618 nsew signal input
rlabel metal2 s 22982 -800 23094 480 8 wbs_dat_i[3]
port 619 nsew signal input
rlabel metal2 s 27710 -800 27822 480 8 wbs_dat_i[4]
port 620 nsew signal input
rlabel metal2 s 31256 -800 31368 480 8 wbs_dat_i[5]
port 621 nsew signal input
rlabel metal2 s 34802 -800 34914 480 8 wbs_dat_i[6]
port 622 nsew signal input
rlabel metal2 s 38348 -800 38460 480 8 wbs_dat_i[7]
port 623 nsew signal input
rlabel metal2 s 41894 -800 42006 480 8 wbs_dat_i[8]
port 624 nsew signal input
rlabel metal2 s 45440 -800 45552 480 8 wbs_dat_i[9]
port 625 nsew signal input
rlabel metal2 s 9980 -800 10092 480 8 wbs_dat_o[0]
port 626 nsew signal output
rlabel metal2 s 50168 -800 50280 480 8 wbs_dat_o[10]
port 627 nsew signal output
rlabel metal2 s 53714 -800 53826 480 8 wbs_dat_o[11]
port 628 nsew signal output
rlabel metal2 s 57260 -800 57372 480 8 wbs_dat_o[12]
port 629 nsew signal output
rlabel metal2 s 60806 -800 60918 480 8 wbs_dat_o[13]
port 630 nsew signal output
rlabel metal2 s 64352 -800 64464 480 8 wbs_dat_o[14]
port 631 nsew signal output
rlabel metal2 s 67898 -800 68010 480 8 wbs_dat_o[15]
port 632 nsew signal output
rlabel metal2 s 71444 -800 71556 480 8 wbs_dat_o[16]
port 633 nsew signal output
rlabel metal2 s 74990 -800 75102 480 8 wbs_dat_o[17]
port 634 nsew signal output
rlabel metal2 s 78536 -800 78648 480 8 wbs_dat_o[18]
port 635 nsew signal output
rlabel metal2 s 82082 -800 82194 480 8 wbs_dat_o[19]
port 636 nsew signal output
rlabel metal2 s 14708 -800 14820 480 8 wbs_dat_o[1]
port 637 nsew signal output
rlabel metal2 s 85628 -800 85740 480 8 wbs_dat_o[20]
port 638 nsew signal output
rlabel metal2 s 89174 -800 89286 480 8 wbs_dat_o[21]
port 639 nsew signal output
rlabel metal2 s 92720 -800 92832 480 8 wbs_dat_o[22]
port 640 nsew signal output
rlabel metal2 s 96266 -800 96378 480 8 wbs_dat_o[23]
port 641 nsew signal output
rlabel metal2 s 99812 -800 99924 480 8 wbs_dat_o[24]
port 642 nsew signal output
rlabel metal2 s 103358 -800 103470 480 8 wbs_dat_o[25]
port 643 nsew signal output
rlabel metal2 s 106904 -800 107016 480 8 wbs_dat_o[26]
port 644 nsew signal output
rlabel metal2 s 110450 -800 110562 480 8 wbs_dat_o[27]
port 645 nsew signal output
rlabel metal2 s 113996 -800 114108 480 8 wbs_dat_o[28]
port 646 nsew signal output
rlabel metal2 s 117542 -800 117654 480 8 wbs_dat_o[29]
port 647 nsew signal output
rlabel metal2 s 19436 -800 19548 480 8 wbs_dat_o[2]
port 648 nsew signal output
rlabel metal2 s 121088 -800 121200 480 8 wbs_dat_o[30]
port 649 nsew signal output
rlabel metal2 s 124634 -800 124746 480 8 wbs_dat_o[31]
port 650 nsew signal output
rlabel metal2 s 24164 -800 24276 480 8 wbs_dat_o[3]
port 651 nsew signal output
rlabel metal2 s 28892 -800 29004 480 8 wbs_dat_o[4]
port 652 nsew signal output
rlabel metal2 s 32438 -800 32550 480 8 wbs_dat_o[5]
port 653 nsew signal output
rlabel metal2 s 35984 -800 36096 480 8 wbs_dat_o[6]
port 654 nsew signal output
rlabel metal2 s 39530 -800 39642 480 8 wbs_dat_o[7]
port 655 nsew signal output
rlabel metal2 s 43076 -800 43188 480 8 wbs_dat_o[8]
port 656 nsew signal output
rlabel metal2 s 46622 -800 46734 480 8 wbs_dat_o[9]
port 657 nsew signal output
rlabel metal2 s 11162 -800 11274 480 8 wbs_sel_i[0]
port 658 nsew signal input
rlabel metal2 s 15890 -800 16002 480 8 wbs_sel_i[1]
port 659 nsew signal input
rlabel metal2 s 20618 -800 20730 480 8 wbs_sel_i[2]
port 660 nsew signal input
rlabel metal2 s 25346 -800 25458 480 8 wbs_sel_i[3]
port 661 nsew signal input
rlabel metal2 s 5252 -800 5364 480 8 wbs_stb_i
port 662 nsew signal input
rlabel metal2 s 6434 -800 6546 480 8 wbs_we_i
port 663 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16016934
string GDS_FILE /home/jona/Desktop/Proyecto_Final/caravan/openlane/user_analog_project_wrapper/runs/24_05_08_11_10/results/signoff/user_analog_project_wrapper.magic.gds
string GDS_START 14765678
<< end >>

