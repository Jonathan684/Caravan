MACRO sky130_fd_pr__pfet_01v8_53Y4NB
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pfet_01v8_53Y4NB ;
  ORIGIN 0.965 5.180 ;
  SIZE 1.930 BY 10.360 ;
  PIN a_n50_n967#
    ANTENNAGATEAREA 5.146700 ;
    ANTENNADIFFAREA 16.343800 ;
    PORT
      LAYER nwell ;
        RECT -1.230 0.625 1.230 5.445 ;
        RECT -1.495 -5.445 1.230 0.625 ;
        RECT -1.495 -10.265 0.965 -5.445 ;
      LAYER li1 ;
        RECT -1.050 5.095 1.050 5.265 ;
        RECT -1.050 0.445 -0.880 5.095 ;
        RECT -0.480 0.445 -0.310 3.085 ;
        RECT 0.310 0.445 0.480 3.085 ;
        RECT -1.315 0.275 0.785 0.445 ;
        RECT -1.315 -9.915 -1.145 0.275 ;
        RECT -1.050 -5.095 -0.880 0.275 ;
        RECT -0.480 -0.065 -0.310 0.275 ;
        RECT -0.515 -0.235 -0.015 -0.065 ;
        RECT -0.745 -5.095 -0.575 -0.450 ;
        RECT -0.480 -3.085 -0.310 -0.235 ;
        RECT 0.045 -4.585 0.215 -0.450 ;
        RECT 0.310 -3.085 0.480 0.275 ;
        RECT -0.250 -4.755 0.250 -4.585 ;
        RECT 0.045 -5.095 0.215 -4.755 ;
        RECT 0.615 -5.095 0.785 0.275 ;
        RECT 0.880 -5.095 1.050 5.095 ;
        RECT -1.050 -5.265 1.050 -5.095 ;
        RECT -0.745 -9.190 -0.575 -5.265 ;
        RECT 0.045 -9.190 0.215 -5.265 ;
        RECT -0.515 -9.575 -0.015 -9.405 ;
        RECT 0.615 -9.915 0.785 -5.265 ;
        RECT -1.315 -10.085 0.785 -9.915 ;
      LAYER met1 ;
        RECT -0.630 5.065 0.630 5.295 ;
        RECT -0.510 -0.035 -0.280 3.065 ;
        RECT 0.280 1.000 0.510 3.065 ;
        RECT 0.000 0.000 1.000 1.000 ;
        RECT -0.510 -0.265 -0.035 -0.035 ;
        RECT -0.775 -9.170 -0.545 -0.470 ;
        RECT -0.510 -3.065 -0.280 -0.265 ;
        RECT 0.015 -1.000 0.245 -0.470 ;
        RECT 0.280 -1.000 0.510 0.000 ;
        RECT 0.000 -2.000 1.000 -1.000 ;
        RECT 0.015 -3.000 0.245 -2.000 ;
        RECT 0.280 -3.000 0.510 -2.000 ;
        RECT 0.000 -4.000 1.000 -3.000 ;
        RECT 0.015 -4.555 0.245 -4.000 ;
        RECT -0.195 -4.785 0.245 -4.555 ;
        RECT 0.015 -5.000 0.245 -4.785 ;
        RECT 0.000 -6.000 1.000 -5.000 ;
        RECT 0.015 -7.000 0.245 -6.000 ;
        RECT 0.000 -8.000 1.000 -7.000 ;
        RECT 0.015 -9.000 0.245 -8.000 ;
        RECT -0.495 -9.605 -0.035 -9.375 ;
        RECT 0.000 -10.000 1.000 -9.000 ;
    END
  END a_n50_n967#
  OBS
      LAYER li1 ;
        RECT -0.250 4.585 0.250 4.755 ;
      LAYER met1 ;
        RECT -0.195 4.555 0.195 4.785 ;
  END
END sky130_fd_pr__pfet_01v8_53Y4NB
END LIBRARY

