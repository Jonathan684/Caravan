VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO inverter
  CLASS BLOCK ;
  FOREIGN inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.670 BY 11.770 ;
  PIN in
    ANTENNAGATEAREA 1.350000 ;
    PORT
      LAYER li1 ;
        RECT 4.930 6.030 5.260 6.200 ;
        RECT 4.450 4.390 4.780 4.560 ;
        RECT 5.410 4.390 5.740 4.560 ;
        RECT 4.975 0.785 5.305 0.955 ;
        RECT 4.495 -1.265 4.825 -1.095 ;
        RECT 5.455 -1.265 5.785 -1.095 ;
      LAYER met1 ;
        RECT 4.950 6.200 5.240 6.230 ;
        RECT 1.840 6.195 5.240 6.200 ;
        RECT 1.795 6.030 5.240 6.195 ;
        RECT 1.795 4.570 2.005 6.030 ;
        RECT 4.950 6.000 5.240 6.030 ;
        RECT 4.470 4.570 4.760 4.590 ;
        RECT 5.430 4.570 5.720 4.590 ;
        RECT 1.795 4.370 5.720 4.570 ;
        RECT 0.000 2.675 1.000 3.180 ;
        RECT 1.795 2.675 2.005 4.370 ;
        RECT 4.470 4.360 4.760 4.370 ;
        RECT 5.430 4.360 5.720 4.370 ;
        RECT 0.000 2.465 2.005 2.675 ;
        RECT 0.000 2.180 1.000 2.465 ;
        RECT 1.795 0.980 2.005 2.465 ;
        RECT 4.995 0.980 5.285 0.985 ;
        RECT 1.795 0.760 5.285 0.980 ;
        RECT 1.795 -1.080 2.005 0.760 ;
        RECT 4.995 0.755 5.285 0.760 ;
        RECT 4.515 -1.080 4.805 -1.065 ;
        RECT 5.475 -1.080 5.765 -1.065 ;
        RECT 1.795 -1.290 5.765 -1.080 ;
        RECT 4.515 -1.295 4.805 -1.290 ;
        RECT 5.475 -1.295 5.765 -1.290 ;
    END
  END in
  PIN gnd
    ANTENNADIFFAREA 2.813500 ;
    PORT
      LAYER pwell ;
        RECT 3.585 -1.955 6.695 1.645 ;
      LAYER li1 ;
        RECT 3.765 1.295 6.515 1.465 ;
        RECT 3.765 -1.605 3.935 1.295 ;
        RECT 4.815 -0.925 4.985 0.615 ;
        RECT 5.775 -0.925 5.945 0.615 ;
        RECT 6.345 -1.605 6.515 1.295 ;
        RECT 3.765 -1.775 6.515 -1.605 ;
      LAYER met1 ;
        RECT 4.785 -0.510 5.015 -0.150 ;
        RECT 5.745 -0.510 5.975 -0.150 ;
        RECT 4.785 -0.760 7.630 -0.510 ;
        RECT 4.785 -0.820 5.015 -0.760 ;
        RECT 5.745 -0.820 5.975 -0.760 ;
        RECT 4.115 -1.580 6.165 -1.575 ;
        RECT 7.350 -1.580 7.620 -0.760 ;
        RECT 2.220 -2.860 7.950 -1.580 ;
        RECT 4.670 -3.470 5.670 -2.860 ;
    END
  END gnd
  PIN Vdd
    ANTENNADIFFAREA 2.376150 ;
    PORT
      LAYER nwell ;
        RECT 3.540 3.700 6.650 6.890 ;
      LAYER li1 ;
        RECT 3.720 6.540 6.470 6.710 ;
        RECT 3.720 4.050 3.890 6.540 ;
        RECT 4.770 4.820 4.940 5.770 ;
        RECT 5.730 4.820 5.900 5.770 ;
        RECT 6.300 4.050 6.470 6.540 ;
        RECT 3.720 3.880 6.470 4.050 ;
      LAYER met1 ;
        RECT 4.440 7.510 5.440 8.300 ;
        RECT 2.500 6.510 7.810 7.510 ;
        RECT 7.140 5.930 7.280 6.510 ;
        RECT 7.130 5.710 7.280 5.930 ;
        RECT 4.710 5.550 7.290 5.710 ;
        RECT 4.740 5.240 4.970 5.550 ;
        RECT 5.700 5.240 5.930 5.550 ;
    END
  END Vdd
  PIN out
    ANTENNADIFFAREA 1.487050 ;
    PORT
      LAYER li1 ;
        RECT 4.290 4.820 4.460 5.770 ;
        RECT 5.250 4.820 5.420 5.770 ;
        RECT 4.335 -0.925 4.505 0.615 ;
        RECT 5.295 -0.925 5.465 0.615 ;
      LAYER met1 ;
        RECT 4.260 5.090 4.490 5.350 ;
        RECT 5.220 5.090 5.450 5.350 ;
        RECT 7.640 5.090 7.790 5.105 ;
        RECT 4.260 4.940 7.790 5.090 ;
        RECT 4.260 4.880 4.490 4.940 ;
        RECT 5.220 4.880 5.450 4.940 ;
        RECT 7.640 2.560 7.790 4.940 ;
        RECT 8.670 2.560 9.670 3.030 ;
        RECT 7.640 2.360 9.670 2.560 ;
        RECT 4.305 0.400 4.535 0.510 ;
        RECT 5.265 0.400 5.495 0.510 ;
        RECT 7.640 0.400 7.790 2.360 ;
        RECT 8.670 2.030 9.670 2.360 ;
        RECT 4.305 0.190 7.800 0.400 ;
        RECT 4.305 0.170 7.630 0.190 ;
        RECT 4.305 -0.160 4.535 0.170 ;
        RECT 5.265 -0.160 5.495 0.170 ;
    END
  END out
END inverter
END LIBRARY

