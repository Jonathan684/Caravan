MACRO example_por
  CLASS BLOCK ;
  FOREIGN example_por ;
  ORIGIN 0.000 0.000 ;
  SIZE 56.720 BY 41.690 ;
  PIN vdd3v3
    ANTENNADIFFAREA 42.573048 ;
    PORT
      LAYER met4 ;
        RECT 0.190 39.825 0.365 41.415 ;
    END
  END vdd3v3
  PIN vdd1v8
    ANTENNADIFFAREA 7.828500 ;
    PORT
      LAYER met4 ;
        RECT 54.870 39.810 55.900 41.455 ;
    END
  END vdd1v8
  PIN vss
    ANTENNADIFFAREA 58.444324 ;
    PORT
      LAYER met4 ;
        RECT 0.190 36.275 1.160 38.275 ;
    END
  END vss
  PIN porb_h
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met3 ;
        RECT 54.845 33.825 56.710 34.170 ;
    END
  END porb_h
  PIN por_l
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met3 ;
        RECT 55.945 37.455 56.720 37.755 ;
    END
  END por_l
  PIN porb_l
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER met3 ;
        RECT 55.940 39.280 56.715 39.580 ;
    END
  END porb_l
  OBS
      LAYER pwell ;
        RECT 0.050 30.500 54.410 30.930 ;
        RECT 0.050 0.480 0.480 30.500 ;
        RECT 0.050 0.050 54.410 0.480 ;
      LAYER li1 ;
        RECT 0.175 0.180 54.300 41.440 ;
      LAYER met1 ;
        RECT 0.125 0.055 54.575 41.430 ;
      LAYER met2 ;
        RECT 0.190 30.880 54.590 41.435 ;
      LAYER met3 ;
        RECT 0.190 39.980 55.945 41.415 ;
        RECT 0.190 38.880 55.540 39.980 ;
        RECT 0.190 38.155 55.945 38.880 ;
        RECT 0.190 37.055 55.545 38.155 ;
        RECT 0.190 34.570 55.945 37.055 ;
        RECT 0.190 33.425 54.445 34.570 ;
        RECT 0.190 0.255 55.945 33.425 ;
      LAYER met4 ;
        RECT 0.765 39.425 54.470 41.455 ;
        RECT 0.365 39.410 54.470 39.425 ;
        RECT 0.365 38.675 55.890 39.410 ;
        RECT 1.560 35.875 55.890 38.675 ;
        RECT 0.365 0.255 55.890 35.875 ;
      LAYER met5 ;
        RECT 21.565 0.250 55.855 38.895 ;
  END
END example_por
END LIBRARY

